module mac_top
(cfg , error , read , rst_n , mac_out , enable , in_b , valid , mode , in_a , clk);
input [15:0] in_a;
input [15:0] in_b;
output [15:0] mac_out;
input clk;
input rst_n;
input enable;
input valid;
input read;
input mode;
input cfg;
output error;
DFFRQX4 \b_reg_reg[7] (.D ( n1036 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[7] ));
DFFRQXL \a_reg_reg[5] (.D ( n1017 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[5] ));
DFFRHQX2 \b_reg_reg[2] (.D ( n1031 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[2] ));
DFFRQX1 \c_reg_reg[14] (.D ( n997 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[14] ));
DFFRQX1 \c_reg_reg[5] (.D ( n1006 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[5] ));
DFFRHQX1 \c_reg_reg[13] (.D ( n998 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[13] ));
ADDFX2 \intadd_7/U4   (.A ( \intadd_7/A[0] ) , .B ( \intadd_7/B[0] ) , .CI ( \intadd_7/CI  ) , .CO ( \intadd_7/n3  ) , .S ( \intadd_7/SUM[0] ));
DFFRX1 \b_reg_reg[6] (.D ( n1035 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[6] ) , .QN ( n2761 ));
DFFRX1 \a_reg_reg[3] (.D ( n1015 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[3] ) , .QN ( n2760 ));
DFFRQX2 \c_reg_reg[1] (.D ( n1010 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[1] ));
DFFRQX2 \c_reg_reg[10] (.D ( n1001 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[10] ));
DFFRQX2 \c_reg_reg[8] (.D ( n1003 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[8] ));
DFFRQX2 \a_reg_reg[6] (.D ( n1018 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[6] ));
DFFRQX1 \c_reg_reg[3] (.D ( n1008 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[3] ));
DFFRQX2 \c_reg_reg[7] (.D ( n1004 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[7] ));
DFFRQX1 \a_reg_reg[14] (.D ( n1026 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[14] ));
DFFRQX1 \b_reg_reg[15] (.D ( n1044 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[15] ));
DFFRQX2 \c_reg_reg[6] (.D ( n1005 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[6] ));
DFFRQX2 \c_reg_reg[0] (.D ( n1011 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[0] ));
DFFRQX2 \c_reg_reg[11] (.D ( n1000 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[11] ));
DFFRQX1 \a_reg_reg[10] (.D ( n1022 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[10] ));
DFFRQX1 \b_reg_reg[10] (.D ( n1039 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[10] ));
DFFRQX1 \b_reg_reg[13] (.D ( n1042 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[13] ));
DFFRQX1 \b_reg_reg[11] (.D ( n1040 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[11] ));
DFFRQX1 \a_reg_reg[13] (.D ( n1025 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[13] ));
DFFRQX1 \a_reg_reg[11] (.D ( n1023 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[11] ));
DFFRQX1 \b_reg_reg[14] (.D ( n1043 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[14] ));
DFFRQX1 \b_reg_reg[12] (.D ( n1041 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[12] ));
DFFRQX1 \a_reg_reg[12] (.D ( n1024 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[12] ));
DFFRQX1 \a_reg_reg[15] (.D ( n1027 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[15] ));
DFFRQX1 \c_reg_reg[15] (.D ( n996 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[15] ));
DFFRQX1 \b_reg_reg[9] (.D ( n1038 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[9] ));
DFFRQX2 \b_reg_reg[5] (.D ( n1034 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[5] ));
DFFRQX2 \b_reg_reg[4] (.D ( n1033 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[4] ));
DFFRHQX4 mode_reg_reg  (.D ( n1028 ) , .CK ( clk ) , .RN ( clk ) , .Q ( \u_mac/mul/multiplier_input2[10] ));
DFFRQX1 \a_reg_reg[8] (.D ( n1020 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[8] ));
DFFRHQX2 \a_reg_reg[2] (.D ( n1014 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[2] ));
DFFRHQX4 \b_reg_reg[0] (.D ( n1029 ) , .CK ( clk ) , .RN ( clk ) , .Q ( \u_mac/mul/N17  ));
DFFRHQX4 \a_reg_reg[0] (.D ( n1012 ) , .CK ( clk ) , .RN ( clk ) , .Q ( \u_mac/mul/N7  ));
DFFRQX1 \c_reg_reg[4] (.D ( n1007 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[4] ));
DFFRQX2 \c_reg_reg[2] (.D ( n1009 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[2] ));
DFFRQX2 \a_reg_reg[9] (.D ( n1021 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[9] ));
DFFRHQX4 \b_reg_reg[1] (.D ( n1030 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[1] ));
DFFRQX2 \c_reg_reg[12] (.D ( n999 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[12] ));
DFFRHQX4 \a_reg_reg[7] (.D ( n1019 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[7] ));
DFFRQX1 \b_reg_reg[8] (.D ( n1037 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[8] ));
ADDFX1 \intadd_4/U4   (.A ( a[12] ) , .B ( b[12] ) , .CI ( \intadd_4/n4  ) , .CO ( \intadd_4/n3  ) , .S ( \intadd_4/SUM[1] ));
ADDFX2 \intadd_7/U3   (.A ( \intadd_7/A[1] ) , .B ( \intadd_7/B[1] ) , .CI ( \intadd_7/n3  ) , .CO ( \intadd_7/n2  ) , .S ( \intadd_7/SUM[1] ));
DFFRHQX4 \a_reg_reg[1] (.D ( n1013 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[1] ));
DFFRQX4 \b_reg_reg[3] (.D ( n1032 ) , .CK ( clk ) , .RN ( clk ) , .Q ( b[3] ));
DFFRQX2 \a_reg_reg[4] (.D ( n1016 ) , .CK ( clk ) , .RN ( clk ) , .Q ( a[4] ));
ADDFX1 \intadd_4/U5   (.A ( a[11] ) , .B ( b[11] ) , .CI ( \intadd_4/CI  ) , .CO ( \intadd_4/n4  ) , .S ( \intadd_4/SUM[0] ));
ADDFX1 \intadd_4/U3   (.A ( a[13] ) , .B ( b[13] ) , .CI ( \intadd_4/n3  ) , .CO ( \intadd_4/n2  ) , .S ( \intadd_4/SUM[2] ));
DFFRQX2 \c_reg_reg[9] (.D ( n1002 ) , .CK ( clk ) , .RN ( clk ) , .Q ( c[9] ));
MX2X1 U959  (.A ( c[9] ) , .B ( n2746 ) , .S0 ( n2749 ) , .Y ( n1002 ));
OAI2BB1X1 U960  (.A0N ( n1048 ) , .A1N ( n2728 ) , .B0 ( n2622 ) , .Y ( n996 ));
AOI22X2 U961  (.A0 ( n2671 ) , .A1 ( n2665 ) , .B0 ( n2659 ) , .B1 ( n2670 ) , .Y ( n2720 ));
AOI21X2 U962  (.A0 ( n2671 ) , .A1 ( n2670 ) , .B0 ( n2669 ) , .Y ( n2719 ));
AOI211X1 U963  (.A0 ( n2692 ) , .A1 ( n2631 ) , .B0 ( n2630 ) , .C0 ( n2629 ) , .Y ( n2714 ));
OAI22XL U964  (.A0 ( n2674 ) , .A1 ( n2658 ) , .B0 ( n2678 ) , .B1 ( n2657 ) , .Y ( n2581 ));
OAI2BB1X1 U965  (.A0N ( n2305 ) , .A1N ( n2661 ) , .B0 ( n2660 ) , .Y ( n2662 ));
OAI21X1 U966  (.A0 ( n2668 ) , .A1 ( n2687 ) , .B0 ( n2667 ) , .Y ( n2669 ));
XOR2X1 U967  (.A ( n2539 ) , .B ( n2538 ) , .Y ( n2547 ));
NOR2X2 U968  (.A ( n2597 ) , .B ( n2596 ) , .Y ( n2725 ));
NAND3XL U969  (.A ( n2633 ) , .B ( n2644 ) , .C ( n2650 ) , .Y ( n2641 ));
NAND3XL U970  (.A ( n2666 ) , .B ( n2305 ) , .C ( n2665 ) , .Y ( n2667 ));
AOI21X1 U971  (.A0 ( n2666 ) , .A1 ( n2663 ) , .B0 ( n2577 ) , .Y ( n2578 ));
INVX2 U972  (.A ( n2659 ) , .Y ( n2668 ));
INVX2 U973  (.A ( n2657 ) , .Y ( n2670 ));
INVX2 U974  (.A ( n2679 ) , .Y ( n2663 ));
INVX1 U975  (.A ( n2689 ) , .Y ( n2650 ));
NAND2X2 U976  (.A ( n2562 ) , .B ( n2564 ) , .Y ( n2628 ));
NAND2BX4 U977  (.AN ( n2642 ) , .B ( n2473 ) , .Y ( n2474 ));
OAI22X1 U978  (.A0 ( n2687 ) , .A1 ( n2674 ) , .B0 ( n2675 ) , .B1 ( n2657 ) , .Y ( n2577 ));
NOR3XL U979  (.A ( n2562 ) , .B ( n2568 ) , .C ( n2561 ) , .Y ( n2563 ));
AOI22XL U980  (.A0 ( n2496 ) , .A1 ( n2636 ) , .B0 ( n2666 ) , .B1 ( n2644 ) , .Y ( n2497 ));
INVX2 U981  (.A ( n2636 ) , .Y ( n2687 ));
NOR2X2 U982  (.A ( n2684 ) , .B ( n2689 ) , .Y ( n2473 ));
NOR2X4 U983  (.A ( n2562 ) , .B ( n2296 ) , .Y ( n2659 ));
CLKAND2X3 U984  (.A ( clk ) , .B ( clk ) , .Y ( n2749 ));
INVX6 U985  (.A ( n2633 ) , .Y ( n2684 ));
NOR2X4 U986  (.A ( n2562 ) , .B ( n2690 ) , .Y ( n2689 ));
BUFX6 U987  (.A ( n2488 ) , .Y ( n2675 ));
INVX2 U988  (.A ( n2510 ) , .Y ( n2625 ));
NAND2X4 U989  (.A ( n2508 ) , .B ( n2644 ) , .Y ( n2633 ));
CLKAND2X4 U990  (.A ( n2508 ) , .B ( n2683 ) , .Y ( n2583 ));
INVX2 U991  (.A ( n2673 ) , .Y ( n2644 ));
AND3X6 U992  (.A ( n2472 ) , .B ( n2471 ) , .C ( n2470 ) , .Y ( n2562 ));
INVX2 U993  (.A ( n2654 ) , .Y ( n2676 ));
NAND2X2 U994  (.A ( n2467 ) , .B ( n2466 ) , .Y ( n2471 ));
NAND3X2 U995  (.A ( n2588 ) , .B ( n2584 ) , .C ( n2591 ) , .Y ( n2460 ));
CLKXOR2X2 U996  (.A ( n2458 ) , .B ( n2457 ) , .Y ( n2683 ));
NAND2X2 U997  (.A ( n2462 ) , .B ( n2461 ) , .Y ( n2469 ));
CLKXOR2X8 U998  (.A ( n2464 ) , .B ( n2452 ) , .Y ( n2591 ));
NAND3XL U999  (.A ( n2444 ) , .B ( n2305 ) , .C ( n2443 ) , .Y ( n2448 ));
NAND2X2 U1000  (.A ( n2441 ) , .B ( n2442 ) , .Y ( n2462 ));
NAND2X1 U1001  (.A ( n2444 ) , .B ( n2296 ) , .Y ( n2441 ));
AND2X4 U1002  (.A ( n2421 ) , .B ( n2419 ) , .Y ( n2466 ));
NOR2X2 U1003  (.A ( n2440 ) , .B ( n2439 ) , .Y ( n2442 ));
AOI21X1 U1004  (.A0 ( n2369 ) , .A1 ( n2294 ) , .B0 ( n2550 ) , .Y ( n2295 ));
NAND2X2 U1005  (.A ( n2411 ) , .B ( n2410 ) , .Y ( n2415 ));
OR2X2 U1006  (.A ( n2374 ) , .B ( n2376 ) , .Y ( n2367 ));
INVX2 U1007  (.A ( n2371 ) , .Y ( n2368 ));
NAND2BX2 U1008  (.AN ( n2325 ) , .B ( n2327 ) , .Y ( n2357 ));
AND3X2 U1009  (.A ( n2411 ) , .B ( n2285 ) , .C ( n2284 ) , .Y ( n2376 ));
OR2X2 U1010  (.A ( n2478 ) , .B ( n2349 ) , .Y ( n2480 ));
OR2X2 U1011  (.A ( n2440 ) , .B ( n2276 ) , .Y ( n2371 ));
CLKAND2X4 U1012  (.A ( n2307 ) , .B ( n2305 ) , .Y ( n2320 ));
INVX2 U1013  (.A ( n2411 ) , .Y ( n2440 ));
OAI21X1 U1014  (.A0 ( n2332 ) , .A1 ( n2550 ) , .B0 ( n2296 ) , .Y ( n2334 ));
AND3X2 U1015  (.A ( n2192 ) , .B ( n2411 ) , .C ( n2191 ) , .Y ( n2308 ));
NAND3X4 U1016  (.A ( n2207 ) , .B ( n2206 ) , .C ( n2205 ) , .Y ( n2333 ));
INVX2 U1017  (.A ( n2339 ) , .Y ( n2345 ));
NAND2X4 U1018  (.A ( n2218 ) , .B ( n2556 ) , .Y ( n2621 ));
AND2X4 U1019  (.A ( n2251 ) , .B ( n2252 ) , .Y ( n2411 ));
INVX2 U1020  (.A ( n2219 ) , .Y ( n2283 ));
BUFX2 U1021  (.A ( n2203 ) , .Y ( n2278 ));
MXI2X1 U1022  (.A ( n2260 ) , .B ( n2266 ) , .S0 ( n2280 ) , .Y ( n2274 ));
CLKXOR2X4 U1023  (.A ( n2200 ) , .B ( n2199 ) , .Y ( n2234 ));
CLKAND2X4 U1024  (.A ( n2275 ) , .B ( n2229 ) , .Y ( n2286 ));
NAND2X6 U1025  (.A ( n2275 ) , .B ( n2280 ) , .Y ( n2269 ));
MXI2X1 U1026  (.A ( n2243 ) , .B ( n2238 ) , .S0 ( n2277 ) , .Y ( n2208 ));
MXI2X2 U1027  (.A ( n2246 ) , .B ( n2245 ) , .S0 ( n2277 ) , .Y ( n2268 ));
AND2X2 U1028  (.A ( n2233 ) , .B ( n2241 ) , .Y ( n2266 ));
CLKXOR2X4 U1029  (.A ( n2183 ) , .B ( n2185 ) , .Y ( n2199 ));
MXI2X1 U1030  (.A ( c[5] ) , .B ( n2329 ) , .S0 ( n2218 ) , .Y ( n2238 ));
INVX10 U1031  (.A ( n2221 ) , .Y ( n2280 ));
BUFX14 U1032  (.A ( n2189 ) , .Y ( n2218 ));
INVX2 U1033  (.A ( n2568 ) , .Y ( n2549 ));
MXI2X4 U1034  (.A ( n2527 ) , .B ( c[13] ) , .S0 ( n2189 ) , .Y ( n2568 ));
NAND2X4 U1035  (.A ( n2170 ) , .B ( n2184 ) , .Y ( n2183 ));
INVX2 U1036  (.A ( n2172 ) , .Y ( n2170 ));
INVX2 U1037  (.A ( n2184 ) , .Y ( n2171 ));
MXI2X4 U1038  (.A ( n2155 ) , .B ( n2154 ) , .S0 ( n2189 ) , .Y ( n2172 ));
MXI2X4 U1039  (.A ( n2149 ) , .B ( n2151 ) , .S0 ( n2189 ) , .Y ( n2160 ));
INVX2 U1040  (.A ( n2163 ) , .Y ( n2162 ));
AND2X2 U1041  (.A ( n2445 ) , .B ( c[10] ) , .Y ( n2163 ));
NOR2X2 U1042  (.A ( n2540 ) , .B ( n2445 ) , .Y ( n2151 ));
CLKNAND2X2 U1043  (.A ( n2139 ) , .B ( n2181 ) , .Y ( n1985 ));
CLKNAND2X8 U1044  (.A ( n2554 ) , .B ( n1984 ) , .Y ( n2181 ));
INVX2 U1045  (.A ( n2187 ) , .Y ( n2418 ));
NAND2X2 U1046  (.A ( n2152 ) , .B ( n2523 ) , .Y ( n2138 ));
INVX10 U1047  (.A ( n2505 ) , .Y ( n2445 ));
NAND2X6 U1048  (.A ( n1983 ) , .B ( n1982 ) , .Y ( n2554 ));
AOI22XL U1049  (.A0 ( n2109 ) , .A1 ( n2108 ) , .B0 ( n2107 ) , .B1 ( n2106 ) , .Y ( n2125 ));
NAND2X2 U1050  (.A ( n1971 ) , .B ( n1961 ) , .Y ( n1969 ));
AND2X6 U1051  (.A ( n1917 ) , .B ( n1916 ) , .Y ( n2505 ));
OAI21X4 U1052  (.A0 ( n2214 ) , .A1 ( n1972 ) , .B0 ( n2211 ) , .Y ( n1971 ));
INVX1 U1053  (.A ( n1977 ) , .Y ( n1979 ));
AOI21X1 U1054  (.A0 ( n1914 ) , .A1 ( n1946 ) , .B0 ( n1913 ) , .Y ( n1915 ));
INVX2 U1055  (.A ( n1934 ) , .Y ( n1946 ));
CLKXOR2X4 U1056  (.A ( n1993 ) , .B ( n1963 ) , .Y ( n2014 ));
CLKXOR2X4 U1057  (.A ( n1909 ) , .B ( n1908 ) , .Y ( n2017 ));
XOR2X4 U1058  (.A ( n1933 ) , .B ( n1932 ) , .Y ( n2213 ));
INVX5 U1059  (.A ( n1888 ) , .Y ( n1993 ));
CLKAND2X3 U1060  (.A ( n1853 ) , .B ( n1854 ) , .Y ( n1895 ));
NAND2X4 U1061  (.A ( n2081 ) , .B ( n2086 ) , .Y ( n1852 ));
CLKNAND2X2 U1062  (.A ( n2055 ) , .B ( n1891 ) , .Y ( n1777 ));
ADDFX1 U1063  (.A ( a[14] ) , .B ( b[14] ) , .CI ( \intadd_4/n2  ) , .CO ( \intadd_4/n1  ) , .S ( \intadd_4/SUM[3] ));
OR2X4 U1064  (.A ( n1806 ) , .B ( n1792 ) , .Y ( n1859 ));
NAND2X5 U1065  (.A ( n1992 ) , .B ( n1996 ) , .Y ( n1889 ));
OAI2BB1X1 U1066  (.A0N ( n1727 ) , .A1N ( n1726 ) , .B0 ( n1767 ) , .Y ( n1771 ));
CLKINVX2 U1067  (.A ( n1805 ) , .Y ( n1792 ));
AOI21X1 U1068  (.A0 ( n1850 ) , .A1 ( n1865 ) , .B0 ( n1849 ) , .Y ( n1862 ));
NAND2X2 U1069  (.A ( n1842 ) , .B ( n1841 ) , .Y ( n1843 ));
CLKAND2X4 U1070  (.A ( n1666 ) , .B ( n1665 ) , .Y ( n1991 ));
INVX1 U1071  (.A ( n1838 ) , .Y ( n1841 ));
INVX2 U1072  (.A ( n1549 ) , .Y ( n1552 ));
NOR2X4 U1073  (.A ( n1548 ) , .B ( n1547 ) , .Y ( n1927 ));
NAND2X2 U1074  (.A ( n1817 ) , .B ( n2702 ) , .Y ( n1838 ));
INVX4 U1075  (.A ( n1672 ) , .Y ( n1673 ));
CLKXOR2X4 U1076  (.A ( n1816 ) , .B ( n1798 ) , .Y ( n1807 ));
NAND2X2 U1077  (.A ( n1743 ) , .B ( n1742 ) , .Y ( n1781 ));
NAND2X2 U1078  (.A ( n1447 ) , .B ( n1446 ) , .Y ( n1907 ));
AOI21X2 U1079  (.A0 ( n1691 ) , .A1 ( n1690 ) , .B0 ( n1694 ) , .Y ( n1730 ));
XOR2X1 U1080  (.A ( n1832 ) , .B ( n1787 ) , .Y ( n1788 ));
NAND3X2 U1081  (.A ( n1816 ) , .B ( n1815 ) , .C ( n1814 ) , .Y ( n1817 ));
CLKNAND2X8 U1082  (.A ( n1769 ) , .B ( n1825 ) , .Y ( n1811 ));
XOR2X1 U1083  (.A ( n1785 ) , .B ( n1752 ) , .Y ( n1779 ));
OAI21X1 U1084  (.A0 ( n1749 ) , .A1 ( n1748 ) , .B0 ( n1747 ) , .Y ( n1785 ));
INVX2 U1085  (.A ( n1641 ) , .Y ( n1644 ));
NOR2X2 U1086  (.A ( n1802 ) , .B ( n1800 ) , .Y ( n1825 ));
XOR2X1 U1087  (.A ( n1681 ) , .B ( n1640 ) , .Y ( n1642 ));
INVX1 U1088  (.A ( n1481 ) , .Y ( n1479 ));
XOR2X1 U1089  (.A ( n1689 ) , .B ( n1745 ) , .Y ( n1741 ));
OAI21X1 U1090  (.A0 ( n1830 ) , .A1 ( n1802 ) , .B0 ( n1688 ) , .Y ( n1745 ));
OAI21X1 U1091  (.A0 ( n1574 ) , .A1 ( n1530 ) , .B0 ( n1621 ) , .Y ( n1532 ));
OAI21X1 U1092  (.A0 ( n1760 ) , .A1 ( n1759 ) , .B0 ( n1758 ) , .Y ( n1794 ));
OAI21X1 U1093  (.A0 ( n1660 ) , .A1 ( a[4] ) , .B0 ( n1760 ) , .Y ( n1720 ));
OAI21X1 U1094  (.A0 ( n1631 ) , .A1 ( n1630 ) , .B0 ( n1629 ) , .Y ( n1679 ));
XOR2X1 U1095  (.A ( n1763 ) , .B ( n1762 ) , .Y ( n1793 ));
NAND2X2 U1096  (.A ( n1835 ) , .B ( n2731 ) , .Y ( n1830 ));
NAND2X2 U1097  (.A ( n1439 ) , .B ( n1440 ) , .Y ( n1418 ));
AOI21X1 U1098  (.A0 ( n1654 ) , .A1 ( n1653 ) , .B0 ( n1652 ) , .Y ( n1721 ));
NAND3XL U1099  (.A ( n1761 ) , .B ( n1818 ) , .C ( n2702 ) , .Y ( n1762 ));
INVX1 U1100  (.A ( n1437 ) , .Y ( n1417 ));
OAI21X1 U1101  (.A0 ( n1617 ) , .A1 ( n1616 ) , .B0 ( n1618 ) , .Y ( n1695 ));
NAND2X2 U1102  (.A ( n1558 ) , .B ( n1557 ) , .Y ( n1569 ));
OAI21X1 U1103  (.A0 ( n1812 ) , .A1 ( n1718 ) , .B0 ( n1717 ) , .Y ( n1756 ));
OA21X1 U1104  (.A0 ( n1656 ) , .A1 ( n1800 ) , .B0 ( n1591 ) , .Y ( n1648 ));
INVX2 U1105  (.A ( n1621 ) , .Y ( n1624 ));
NAND2X2 U1106  (.A ( n1635 ) , .B ( n1636 ) , .Y ( n1748 ));
NAND2X2 U1107  (.A ( n1660 ) , .B ( a[4] ) , .Y ( n1760 ));
AOI21X4 U1108  (.A0 ( n1400 ) , .A1 ( n1409 ) , .B0 ( n1407 ) , .Y ( n1449 ));
NAND3X2 U1109  (.A ( n1711 ) , .B ( n1710 ) , .C ( n1714 ) , .Y ( n1763 ));
AND2X2 U1110  (.A ( n1659 ) , .B ( n1658 ) , .Y ( n1660 ));
OAI21X1 U1111  (.A0 ( n1599 ) , .A1 ( n1118 ) , .B0 ( n1598 ) , .Y ( n1652 ));
OAI21X1 U1112  (.A0 ( n1594 ) , .A1 ( n1593 ) , .B0 ( n1592 ) , .Y ( n1595 ));
AOI21XL U1113  (.A0 ( n2703 ) , .A1 ( n2706 ) , .B0 ( n2707 ) , .Y ( \intadd_7/B[2] ));
OAI21XL U1114  (.A0 ( n1656 ) , .A1 ( n1655 ) , .B0 ( n1761 ) , .Y ( n1659 ));
XOR2X1 U1115  (.A ( n1634 ) , .B ( n1633 ) , .Y ( n1635 ));
INVX2 U1116  (.A ( n1819 ) , .Y ( n1802 ));
AOI21X2 U1117  (.A0 ( n1467 ) , .A1 ( n1466 ) , .B0 ( n1465 ) , .Y ( n1469 ));
CLKXOR2X2 U1118  (.A ( n1599 ) , .B ( n1543 ) , .Y ( n1594 ));
CLKXOR2X4 U1119  (.A ( n1194 ) , .B ( n1193 ) , .Y ( n1195 ));
NAND3X2 U1120  (.A ( n1380 ) , .B ( n1379 ) , .C ( n1378 ) , .Y ( n1381 ));
NAND2X2 U1121  (.A ( n1424 ) , .B ( n2748 ) , .Y ( n1539 ));
CLKXOR2X4 U1122  (.A ( n1056 ) , .B ( n1279 ) , .Y ( n1282 ));
XOR2X1 U1123  (.A ( n1340 ) , .B ( n1339 ) , .Y ( n1193 ));
OAI21X1 U1124  (.A0 ( n1118 ) , .A1 ( n1800 ) , .B0 ( n1488 ) , .Y ( n1494 ));
INVX2 U1125  (.A ( n1049 ) , .Y ( n1823 ));
NAND2X5 U1126  (.A ( n1338 ) , .B ( n1340 ) , .Y ( n1374 ));
NAND2X4 U1127  (.A ( n1337 ) , .B ( n1339 ) , .Y ( n1376 ));
XOR2X1 U1128  (.A ( n1078 ) , .B ( n2706 ) , .Y ( n1280 ));
XOR2X1 U1129  (.A ( n2701 ) , .B ( n2700 ) , .Y ( n2704 ));
INVX2 U1130  (.A ( n1818 ) , .Y ( n1655 ));
CLKXOR2X4 U1131  (.A ( n1192 ) , .B ( n1301 ) , .Y ( n1339 ));
AOI21X1 U1132  (.A0 ( n1274 ) , .A1 ( n1273 ) , .B0 ( n1272 ) , .Y ( n1275 ));
NAND2X4 U1133  (.A ( n1199 ) , .B ( n1167 ) , .Y ( n1338 ));
INVX2 U1134  (.A ( n1267 ) , .Y ( n1458 ));
NAND2X5 U1135  (.A ( a[9] ) , .B ( n2293 ) , .Y ( n1049 ));
NOR3X1 U1136  (.A ( n1260 ) , .B ( n1259 ) , .C ( n1686 ) , .Y ( n1261 ));
XOR2X3 U1137  (.A ( n1326 ) , .B ( n1305 ) , .Y ( n1308 ));
CLKAND2X4 U1138  (.A ( n1464 ) , .B ( n1322 ) , .Y ( n1327 ));
INVX4 U1139  (.A ( n1800 ) , .Y ( n1820 ));
XOR2X1 U1140  (.A ( n1269 ) , .B ( n1101 ) , .Y ( n1102 ));
NAND2BX2 U1141  (.AN ( n1181 ) , .B ( n1179 ) , .Y ( n1302 ));
CLKAND2X4 U1142  (.A ( n1326 ) , .B ( n1191 ) , .Y ( n1301 ));
NAND2X4 U1143  (.A ( b[8] ) , .B ( n2293 ) , .Y ( n1800 ));
NAND2BX4 U1144  (.AN ( n1189 ) , .B ( n1188 ) , .Y ( n1326 ));
NAND2X6 U1145  (.A ( n1144 ) , .B ( n1143 ) , .Y ( n1159 ));
NOR2X2 U1146  (.A ( n1091 ) , .B ( n1487 ) , .Y ( n1098 ));
CLKXOR2X4 U1147  (.A ( n1187 ) , .B ( n1186 ) , .Y ( n1188 ));
INVX2 U1148  (.A ( n2732 ) , .Y ( n1706 ));
INVX2 U1149  (.A ( n1160 ) , .Y ( n1142 ));
CLKXOR2X4 U1150  (.A ( n1070 ) , .B ( n1633 ) , .Y ( n2699 ));
INVX2 U1151  (.A ( b[4] ) , .Y ( n1633 ));
NAND2X2 U1152  (.A ( n1062 ) , .B ( n1061 ) , .Y ( n1877 ));
INVX2 U1153  (.A ( b[5] ) , .Y ( n1061 ));
INVX2 U1154  (.A ( a[6] ) , .Y ( n1075 ));
NAND2BX4 U1155  (.AN ( n1074 ) , .B ( n1759 ) , .Y ( n1882 ));
CLKNAND2X4 U1156  (.A ( n1095 ) , .B ( n1093 ) , .Y ( n1072 ));
INVX4 U1157  (.A ( n1095 ) , .Y ( n1066 ));
INVX2 U1158  (.A ( b[2] ) , .Y ( n1580 ));
NAND2BX2 U1159  (.AN ( n1119 ) , .B ( n1112 ) , .Y ( n1113 ));
BUFX5 U1160  (.A ( \u_mac/mul/N7  ) , .Y ( n2748 ));
XOR2X3 U1161  (.A ( n1089 ) , .B ( a[1] ) , .Y ( n1090 ));
CLKXOR2X2 U1162  (.A ( n1086 ) , .B ( n1085 ) , .Y ( n1087 ));
INVX8 U1163  (.A ( n1119 ) , .Y ( n1107 ));
BUFX8 U1164  (.A ( \u_mac/mul/N17  ) , .Y ( n2750 ));
INVX8 U1165  (.A ( \u_mac/mul/multiplier_input2[10] ) , .Y ( n2643 ));
INVXL U1166  (.A ( n1118 ) , .Y ( n1264 ));
NAND2BX2 U1167  (.AN ( n1118 ) , .B ( n2731 ) , .Y ( n1456 ));
NOR2XL U1168  (.A ( n2697 ) , .B ( n1353 ) , .Y ( n1078 ));
INVXL U1169  (.A ( n1328 ) , .Y ( n1329 ));
INVXL U1170  (.A ( n2706 ) , .Y ( n2708 ));
NOR2XL U1171  (.A ( n2751 ) , .B ( n2735 ) , .Y ( \intadd_7/CI  ));
INVXL U1172  (.A ( \intadd_7/SUM[2] ) , .Y ( n1557 ));
NOR2XL U1173  (.A ( n1288 ) , .B ( n2697 ) , .Y ( n2696 ));
NAND2BXL U1174  (.AN ( n1525 ) , .B ( n1524 ) , .Y ( n1526 ));
INVXL U1175  (.A ( n1528 ) , .Y ( n1578 ));
NAND2XL U1176  (.A ( n2733 ) , .B ( n1657 ) , .Y ( n1705 ));
OAI21X1 U1177  (.A0 ( n1618 ) , .A1 ( n1617 ) , .B0 ( n1695 ) , .Y ( n1678 ));
INVXL U1178  (.A ( n1179 ) , .Y ( n1180 ));
INVXL U1179  (.A ( n1377 ) , .Y ( n1378 ));
NAND2BXL U1180  (.AN ( n1685 ) , .B ( b[4] ) , .Y ( n1751 ));
INVXL U1181  (.A ( n1541 ) , .Y ( n1542 ));
NAND2XL U1182  (.A ( n1250 ) , .B ( n2293 ) , .Y ( n1251 ));
INVXL U1183  (.A ( n1751 ) , .Y ( n1784 ));
OR3XL U1184  (.A ( n1542 ) , .B ( n1118 ) , .C ( n1655 ) , .Y ( n1543 ));
NAND2XL U1185  (.A ( n1811 ) , .B ( n1810 ) , .Y ( n1808 ));
NAND2X4 U1186  (.A ( n2643 ) , .B ( a[7] ) , .Y ( n1088 ));
INVX2 U1187  (.A ( n1176 ) , .Y ( n2732 ));
NAND2XL U1188  (.A ( n1828 ) , .B ( n1845 ) , .Y ( n1839 ));
NOR2X4 U1189  (.A ( n1403 ) , .B ( n1119 ) , .Y ( n1120 ));
INVXL U1190  (.A ( n1214 ) , .Y ( n1217 ));
INVXL U1191  (.A ( n2165 ) , .Y ( n2167 ));
NAND2XL U1192  (.A ( n1539 ) , .B ( n1426 ) , .Y ( n1445 ));
AND2X4 U1193  (.A ( n2160 ) , .B ( n2159 ) , .Y ( n2168 ));
NAND2XL U1194  (.A ( n1388 ) , .B ( n1389 ) , .Y ( n1222 ));
AND2X4 U1195  (.A ( n1856 ) , .B ( n1855 ) , .Y ( n1900 ));
NAND2BXL U1196  (.AN ( n2239 ) , .B ( n2267 ) , .Y ( n2271 ));
CLKAND2X3 U1197  (.A ( n2147 ) , .B ( n2162 ) , .Y ( n2277 ));
INVXL U1198  (.A ( n2376 ) , .Y ( n2377 ));
INVXL U1199  (.A ( n2297 ) , .Y ( n2294 ));
INVXL U1200  (.A ( n1974 ) , .Y ( n1970 ));
OAI21X1 U1201  (.A0 ( n2137 ) , .A1 ( n2136 ) , .B0 ( n2181 ) , .Y ( n2142 ));
AOI21X1 U1202  (.A0 ( n2327 ) , .A1 ( n2564 ) , .B0 ( n2326 ) , .Y ( n2358 ));
AOI2BB2XL U1203  (.B0 ( c[8] ) , .B1 ( n2692 ) , .A0N ( n2297 ) , .A1N ( n2296 ) , .Y ( n2298 ));
NAND2X2 U1204  (.A ( n2417 ) , .B ( n2416 ) , .Y ( n2421 ));
NOR2XL U1205  (.A ( n2522 ) , .B ( n2556 ) , .Y ( n2525 ));
NAND2XL U1206  (.A ( n2476 ) , .B ( n2475 ) , .Y ( n2477 ));
AOI21X1 U1207  (.A0 ( c[11] ) , .A1 ( n2540 ) , .B0 ( n2520 ) , .Y ( n2521 ));
INVXL U1208  (.A ( n2571 ) , .Y ( n2516 ));
NOR2XL U1209  (.A ( \intadd_4/n1  ) , .B ( n1960 ) , .Y ( n1081 ));
XNOR2X1 U1210  (.A ( n2617 ) , .B ( n2594 ) , .Y ( n2726 ));
NAND2BXL U1211  (.AN ( \intadd_4/SUM[3] ) , .B ( n1081 ) , .Y ( n1082 ));
MX2X1 U1212  (.A ( c[8] ) , .B ( n2747 ) , .S0 ( n2749 ) , .Y ( n1003 ));
CLKBUFX4 U1213  (.A ( n2643 ) , .Y ( n2692 ));
BUFX10 U1214  (.A ( n2293 ) , .Y ( n2556 ));
MXI2X2 U1215  (.A ( n2718 ) , .B ( n2580 ) , .S0 ( n2655 ) , .Y ( n1007 ));
AOI222X4 U1216  (.A0 ( n2671 ) , .A1 ( n2683 ) , .B0 ( n2654 ) , .B1 ( n2659 ) , .C0 ( n2579 ) , .C1 ( n2305 ) , .Y ( n2718 ));
NAND2X5 U1217  (.A ( n2434 ) , .B ( n2433 ) , .Y ( n2436 ));
NAND2X2 U1218  (.A ( n2434 ) , .B ( n2435 ) , .Y ( n2400 ));
NAND2X4 U1219  (.A ( n2397 ) , .B ( n2396 ) , .Y ( n2406 ));
OR3X8 U1220  (.A ( n2374 ) , .B ( n2368 ) , .C ( n2376 ) , .Y ( n2369 ));
INVX2 U1221  (.A ( n2239 ) , .Y ( n2202 ));
INVX2 U1222  (.A ( n2279 ) , .Y ( n2204 ));
XOR2XL U1223  (.A ( n2468 ) , .B ( n2446 ) , .Y ( n2447 ));
OAI21X6 U1224  (.A0 ( n2214 ) , .A1 ( n1956 ) , .B0 ( n2211 ) , .Y ( n1943 ));
CLKINVX2 U1225  (.A ( n2040 ) , .Y ( n2044 ));
NAND2X2 U1226  (.A ( n1996 ) , .B ( n1995 ) , .Y ( n1997 ));
NAND2X4 U1227  (.A ( n1609 ) , .B ( n1672 ) , .Y ( n1646 ));
INVX8 U1228  (.A ( n1606 ) , .Y ( n1670 ));
NAND2X6 U1229  (.A ( n1448 ) , .B ( n1907 ) , .Y ( n1931 ));
NAND2X2 U1230  (.A ( n1907 ) , .B ( n1906 ) , .Y ( n1908 ));
NAND2X4 U1231  (.A ( n1605 ) , .B ( n1736 ) , .Y ( n1669 ));
NAND2X4 U1232  (.A ( n1586 ) , .B ( n1585 ) , .Y ( n1734 ));
NAND2X2 U1233  (.A ( n1439 ) , .B ( n1438 ) , .Y ( n1441 ));
NAND2X4 U1234  (.A ( n1531 ) , .B ( n1532 ) , .Y ( n1605 ));
CLKNAND2X2 U1235  (.A ( n2078 ) , .B ( n2106 ) , .Y ( n2095 ));
NAND2X2 U1236  (.A ( n1563 ) , .B ( n1561 ) , .Y ( n1566 ));
INVX4 U1237  (.A ( n1350 ) , .Y ( n1352 ));
OAI21X4 U1238  (.A0 ( n1769 ) , .A1 ( n1825 ) , .B0 ( n1811 ) , .Y ( n1774 ));
NAND2X4 U1239  (.A ( n1382 ) , .B ( n1381 ) , .Y ( n1383 ));
NAND2X4 U1240  (.A ( n1388 ) , .B ( n1387 ) , .Y ( n1390 ));
NAND2X2 U1241  (.A ( n1370 ) , .B ( n1369 ) , .Y ( n1373 ));
AND2X4 U1242  (.A ( n1223 ) , .B ( n1225 ) , .Y ( n1387 ));
NAND3X2 U1243  (.A ( n1376 ) , .B ( n1375 ) , .C ( n1374 ) , .Y ( n1380 ));
NAND2X4 U1244  (.A ( n1376 ) , .B ( n1374 ) , .Y ( n1370 ));
NAND2X6 U1245  (.A ( n1377 ) , .B ( n1375 ) , .Y ( n1371 ));
NAND2BX2 U1246  (.AN ( n1781 ) , .B ( n1780 ) , .Y ( n1790 ));
XOR2X3 U1247  (.A ( n1201 ) , .B ( n1200 ) , .Y ( n1220 ));
NAND2X1 U1248  (.A ( n1228 ) , .B ( n1227 ) , .Y ( n1230 ));
NAND2X4 U1249  (.A ( n1359 ) , .B ( n1360 ) , .Y ( n1357 ));
INVX4 U1250  (.A ( n1166 ) , .Y ( n1199 ));
NAND2X3 U1251  (.A ( n1332 ) , .B ( n1333 ) , .Y ( n1312 ));
INVX4 U1252  (.A ( n1460 ) , .Y ( n1461 ));
INVX4 U1253  (.A ( n1168 ) , .Y ( n1171 ));
INVX4 U1254  (.A ( n1201 ) , .Y ( n1360 ));
INVX1 U1255  (.A ( n1341 ) , .Y ( n1342 ));
AND2X4 U1256  (.A ( n1354 ) , .B ( n1353 ) , .Y ( n1367 ));
INVX2 U1257  (.A ( n1291 ) , .Y ( n1293 ));
OAI21X2 U1258  (.A0 ( n1523 ) , .A1 ( n1522 ) , .B0 ( n1521 ) , .Y ( n1579 ));
NOR2X4 U1259  (.A ( n1263 ) , .B ( n1262 ) , .Y ( n1291 ));
CLKNAND2X2 U1260  (.A ( n1707 ) , .B ( n1582 ) , .Y ( n1313 ));
OAI21XL U1261  (.A0 ( n2692 ) , .A1 ( n1430 ) , .B0 ( n1425 ) , .Y ( n1426 ));
NAND2X1 U1262  (.A ( n2619 ) , .B ( n2290 ) , .Y ( n2292 ));
CLKAND2X2 U1263  (.A ( n1868 ) , .B ( n1867 ) , .Y ( n2117 ));
INVX2 U1264  (.A ( n2733 ) , .Y ( n1177 ));
INVX1 U1265  (.A ( n1636 ) , .Y ( n1637 ));
XOR2X2 U1266  (.A ( n1125 ) , .B ( n1148 ) , .Y ( n1160 ));
OR2XL U1267  (.A ( n1882 ) , .B ( n1881 ) , .Y ( n1883 ));
CLKNAND2X2 U1268  (.A ( n1867 ) , .B ( n1821 ) , .Y ( n1828 ));
INVX1 U1269  (.A ( n1867 ) , .Y ( n1850 ));
INVX1 U1270  (.A ( n1976 ) , .Y ( n1961 ));
INVX2 U1271  (.A ( n1273 ) , .Y ( n1257 ));
NAND2XL U1272  (.A ( n1582 ) , .B ( n1819 ) , .Y ( n1473 ));
INVX2 U1273  (.A ( n1456 ) , .Y ( n1457 ));
INVX1 U1274  (.A ( n1825 ) , .Y ( n1826 ));
INVX4 U1275  (.A ( n2699 ) , .Y ( n1575 ));
NAND2X1 U1276  (.A ( n1824 ) , .B ( n1823 ) , .Y ( n1827 ));
OR2XL U1277  (.A ( n1877 ) , .B ( n1876 ) , .Y ( n1884 ));
OAI21XL U1278  (.A0 ( n1800 ) , .A1 ( n1049 ) , .B0 ( n1822 ) , .Y ( n1801 ));
CLKNAND2X2 U1279  (.A ( n1819 ) , .B ( n1818 ) , .Y ( n1822 ));
CLKAND2X2 U1280  (.A ( b[1] ) , .B ( n2556 ) , .Y ( n1476 ));
INVX4 U1281  (.A ( n1084 ) , .Y ( n1064 ));
AOI21X4 U1282  (.A0 ( n2502 ) , .A1 ( n2556 ) , .B0 ( n1053 ) , .Y ( n2715 ));
OAI22X2 U1283  (.A0 ( n2652 ) , .A1 ( n2651 ) , .B0 ( n2673 ) , .B1 ( n2650 ) , .Y ( n2653 ));
INVX2 U1284  (.A ( n2623 ) , .Y ( n2624 ));
INVX1 U1285  (.A ( n2675 ) , .Y ( n2490 ));
NAND2X2 U1286  (.A ( n2659 ) , .B ( n2561 ) , .Y ( n2597 ));
INVX4 U1287  (.A ( n2591 ) , .Y ( n2688 ));
AOI21X4 U1288  (.A0 ( n2425 ) , .A1 ( n2423 ) , .B0 ( n2405 ) , .Y ( n2409 ));
NAND2X4 U1289  (.A ( n2428 ) , .B ( n2404 ) , .Y ( n2425 ));
NAND2X4 U1290  (.A ( n2426 ) , .B ( n2485 ) , .Y ( n2458 ));
NAND2X4 U1291  (.A ( n2394 ) , .B ( n2373 ) , .Y ( n2407 ));
NAND2X5 U1292  (.A ( n2354 ) , .B ( n2491 ) , .Y ( n2486 ));
INVX2 U1293  (.A ( n2493 ) , .Y ( n2494 ));
NAND2X4 U1294  (.A ( n2323 ) , .B ( n2322 ) , .Y ( n2485 ));
INVX6 U1295  (.A ( n2369 ) , .Y ( n2287 ));
NAND2X4 U1296  (.A ( n2374 ) , .B ( n2305 ) , .Y ( n2378 ));
NAND4X6 U1297  (.A ( n2333 ) , .B ( n2339 ) , .C ( n2340 ) , .D ( n2317 ) , .Y ( n2307 ));
AND2X6 U1298  (.A ( n2231 ) , .B ( n2230 ) , .Y ( n2339 ));
INVX4 U1299  (.A ( n2251 ) , .Y ( n2235 ));
NAND2X2 U1300  (.A ( n2275 ) , .B ( n2274 ) , .Y ( n2276 ));
XOR2X8 U1301  (.A ( n2169 ) , .B ( n2168 ) , .Y ( n2221 ));
NAND2X4 U1302  (.A ( n2167 ) , .B ( n2166 ) , .Y ( n2169 ));
NAND2X4 U1303  (.A ( n2160 ) , .B ( n2148 ) , .Y ( n2156 ));
NAND2X5 U1304  (.A ( n2543 ) , .B ( n2162 ) , .Y ( n2166 ));
INVX6 U1305  (.A ( n2504 ) , .Y ( n2543 ));
AO21XL U1306  (.A0 ( n2614 ) , .A1 ( n2613 ) , .B0 ( n2612 ) , .Y ( n2615 ));
CLKNAND2X2 U1307  (.A ( n2525 ) , .B ( n2524 ) , .Y ( n2592 ));
INVXL U1308  (.A ( n2300 ) , .Y ( n2301 ));
NAND2X2 U1309  (.A ( n2113 ) , .B ( n2112 ) , .Y ( n2114 ));
INVX4 U1310  (.A ( n1900 ) , .Y ( n2082 ));
INVX2 U1311  (.A ( n1669 ) , .Y ( n1671 ));
OAI21X4 U1312  (.A0 ( n1560 ) , .A1 ( n1567 ) , .B0 ( n1559 ) , .Y ( n1573 ));
NAND2X4 U1313  (.A ( n1864 ) , .B ( n1863 ) , .Y ( n2112 ));
INVX2 U1314  (.A ( n1562 ) , .Y ( n1564 ));
INVX3 U1315  (.A ( n1449 ) , .Y ( n1555 ));
NAND2X4 U1316  (.A ( n1405 ) , .B ( n1404 ) , .Y ( n1402 ));
INVX4 U1317  (.A ( n1568 ) , .Y ( n1563 ));
NAND2X2 U1318  (.A ( n1218 ) , .B ( n1227 ) , .Y ( n1225 ));
CLKXOR2X2 U1319  (.A ( n1584 ) , .B ( n1620 ) , .Y ( n1587 ));
INVX2 U1320  (.A ( n1620 ) , .Y ( n1625 ));
NAND2X4 U1321  (.A ( n1530 ) , .B ( n1574 ) , .Y ( n1621 ));
CLKXOR2X2 U1322  (.A ( n1592 ) , .B ( n1544 ) , .Y ( n1545 ));
NAND2X2 U1323  (.A ( n1306 ) , .B ( n1152 ) , .Y ( n1155 ));
INVXL U1324  (.A ( n2036 ) , .Y ( n1242 ));
INVX1 U1325  (.A ( n1445 ) , .Y ( n1446 ));
INVX4 U1326  (.A ( n1152 ) , .Y ( n1154 ));
AND2X2 U1327  (.A ( n1325 ) , .B ( n1323 ) , .Y ( n1305 ));
CLKNAND2X2 U1328  (.A ( n2698 ) , .B ( n1706 ) , .Y ( n1317 ));
XOR2XL U1329  (.A ( n1539 ) , .B ( n1497 ) , .Y ( n1498 ));
INVX2 U1330  (.A ( n1635 ) , .Y ( n1638 ));
INVX2 U1331  (.A ( n1321 ) , .Y ( n1316 ));
NOR2X2 U1332  (.A ( n1458 ) , .B ( n1456 ) , .Y ( n1278 ));
INVXL U1333  (.A ( n1830 ) , .Y ( n1831 ));
XOR2XL U1334  (.A ( n1518 ) , .B ( n1523 ) , .Y ( n1477 ));
AND2X2 U1335  (.A ( n1423 ) , .B ( n1422 ) , .Y ( n1424 ));
NOR2X1 U1336  (.A ( n1172 ) , .B ( n1148 ) , .Y ( n1149 ));
NAND2X2 U1337  (.A ( n1083 ) , .B ( n1082 ) , .Y ( error ));
INVX1 U1338  (.A ( n1323 ) , .Y ( n1324 ));
INVXL U1339  (.A ( n1433 ) , .Y ( n1434 ));
NAND2X2 U1340  (.A ( n1492 ) , .B ( n1818 ) , .Y ( n1488 ));
INVX1 U1341  (.A ( n1822 ) , .Y ( n1824 ));
NAND2BXL U1342  (.AN ( \intadd_4/SUM[2] ) , .B ( n1958 ) , .Y ( n1959 ));
AND2X2 U1343  (.A ( n1121 ) , .B ( n2702 ) , .Y ( n1323 ));
NAND2X2 U1344  (.A ( n1069 ) , .B ( n1107 ) , .Y ( n1070 ));
NAND2X4 U1345  (.A ( n1108 ) , .B ( n1107 ) , .Y ( n1110 ));
NAND2X4 U1346  (.A ( n1106 ) , .B ( n1109 ) , .Y ( n1069 ));
INVXL U1347  (.A ( n1246 ) , .Y ( n1247 ));
OAI21X2 U1348  (.A0 ( n2687 ) , .A1 ( n2686 ) , .B0 ( n2685 ) , .Y ( n2691 ));
OAI21X2 U1349  (.A0 ( n2686 ) , .A1 ( n2658 ) , .B0 ( n2637 ) , .Y ( n2639 ));
NAND2X2 U1350  (.A ( n2642 ) , .B ( n2675 ) , .Y ( n2539 ));
NAND2X2 U1351  (.A ( n2741 ) , .B ( n2749 ) , .Y ( n2566 ));
NAND2X2 U1352  (.A ( n2565 ) , .B ( n2564 ) , .Y ( n2741 ));
NAND2X2 U1353  (.A ( n2659 ) , .B ( n2683 ) , .Y ( n2660 ));
NOR2X4 U1354  (.A ( n2584 ) , .B ( n2677 ) , .Y ( n2453 ));
NAND2X4 U1355  (.A ( n2437 ) , .B ( n2465 ) , .Y ( n2452 ));
NAND3X4 U1356  (.A ( n2401 ) , .B ( n2428 ) , .C ( n2426 ) , .Y ( n2384 ));
NAND2X2 U1357  (.A ( n2429 ) , .B ( n2428 ) , .Y ( n2430 ));
NAND2X4 U1358  (.A ( n2413 ) , .B ( n2295 ) , .Y ( n2299 ));
NAND2X2 U1359  (.A ( n2485 ) , .B ( n2484 ) , .Y ( n2487 ));
NAND2X4 U1360  (.A ( n2331 ) , .B ( n2359 ) , .Y ( n2428 ));
NAND2X2 U1361  (.A ( n2492 ) , .B ( n2491 ) , .Y ( n2495 ));
INVX2 U1362  (.A ( n2658 ) , .Y ( n2665 ));
NAND2X2 U1363  (.A ( n2480 ) , .B ( n2479 ) , .Y ( n2482 ));
INVX2 U1364  (.A ( n2357 ) , .Y ( n2362 ));
OAI21X4 U1365  (.A0 ( n2374 ) , .A1 ( n2550 ) , .B0 ( n2296 ) , .Y ( n2375 ));
NAND2X4 U1366  (.A ( n2478 ) , .B ( n2349 ) , .Y ( n2479 ));
NOR2X6 U1367  (.A ( n2308 ) , .B ( n2307 ) , .Y ( n2325 ));
NOR2X2 U1368  (.A ( n2360 ) , .B ( n2359 ) , .Y ( n2361 ));
INVX2 U1369  (.A ( n2415 ) , .Y ( n2412 ));
MXI2X2 U1370  (.A ( n2194 ) , .B ( n2439 ) , .S0 ( n2235 ) , .Y ( n2207 ));
NAND2BX2 U1371  (.AN ( n2259 ) , .B ( n2283 ) , .Y ( n2284 ));
XOR2X8 U1372  (.A ( n2180 ) , .B ( n2196 ) , .Y ( n2251 ));
NAND2X4 U1373  (.A ( n2197 ) , .B ( n2195 ) , .Y ( n2180 ));
NAND2X4 U1374  (.A ( n2203 ) , .B ( n2221 ) , .Y ( n2239 ));
NAND2X2 U1375  (.A ( n2280 ) , .B ( n2279 ) , .Y ( n2281 ));
MXI2X2 U1376  (.A ( n2246 ) , .B ( n2237 ) , .S0 ( n2241 ) , .Y ( n2219 ));
MXI2X1 U1377  (.A ( c[9] ) , .B ( n2418 ) , .S0 ( n2621 ) , .Y ( n2420 ));
MXI2X3 U1378  (.A ( n2505 ) , .B ( n2632 ) , .S0 ( n2218 ) , .Y ( n2627 ));
INVX2 U1379  (.A ( n2244 ) , .Y ( n2245 ));
MXI2X2 U1380  (.A ( c[4] ) , .B ( n2313 ) , .S0 ( n2218 ) , .Y ( n2243 ));
MXI2X1 U1381  (.A ( c[3] ) , .B ( n2321 ) , .S0 ( n2218 ) , .Y ( n2242 ));
AND2XL U1382  (.A ( n2610 ) , .B ( n2613 ) , .Y ( n2616 ));
INVXL U1383  (.A ( n2572 ) , .Y ( n2576 ));
NAND2X1 U1384  (.A ( n2558 ) , .B ( n2557 ) , .Y ( n2611 ));
INVXL U1385  (.A ( n2527 ) , .Y ( n2528 ));
NAND2BX4 U1386  (.AN ( n2418 ) , .B ( c[9] ) , .Y ( n2132 ));
INVXL U1387  (.A ( n2554 ) , .Y ( n2555 ));
AND2X2 U1388  (.A ( n2445 ) , .B ( n2540 ) , .Y ( n2157 ));
INVXL U1389  (.A ( n2346 ) , .Y ( n2347 ));
XOR2X2 U1390  (.A ( n2122 ) , .B ( n2121 ) , .Y ( n2123 ));
NAND2X4 U1391  (.A ( n2055 ) , .B ( n2057 ) , .Y ( n1894 ));
AND2X2 U1392  (.A ( n1979 ) , .B ( n1978 ) , .Y ( n1980 ));
NAND2X4 U1393  (.A ( n1861 ) , .B ( n1860 ) , .Y ( n2083 ));
INVX4 U1394  (.A ( n2007 ) , .Y ( n2016 ));
NAND2X4 U1395  (.A ( n1770 ) , .B ( n1771 ) , .Y ( n2042 ));
INVX4 U1396  (.A ( n1853 ) , .Y ( n1856 ));
INVX6 U1397  (.A ( n2213 ) , .Y ( n2018 ));
OAI21X4 U1398  (.A0 ( n1755 ) , .A1 ( n1754 ) , .B0 ( n1806 ) , .Y ( n1776 ));
NAND2X4 U1399  (.A ( n1673 ) , .B ( n1728 ) , .Y ( n1675 ));
XOR2X4 U1400  (.A ( n1670 ) , .B ( n1535 ) , .Y ( n1549 ));
AOI21X4 U1401  (.A0 ( n1732 ) , .A1 ( n1731 ) , .B0 ( n1730 ) , .Y ( n1739 ));
NAND2X4 U1402  (.A ( n1534 ) , .B ( n1533 ) , .Y ( n1733 ));
NAND2X4 U1403  (.A ( n1479 ) , .B ( n1478 ) , .Y ( n1502 ));
INVX4 U1404  (.A ( n1531 ) , .Y ( n1534 ));
INVX4 U1405  (.A ( n2086 ) , .Y ( n2111 ));
NAND2BX8 U1406  (.AN ( n1864 ) , .B ( n1862 ) , .Y ( n2086 ));
NAND2X4 U1407  (.A ( n1449 ) , .B ( n1450 ) , .Y ( n1505 ));
NAND2X2 U1408  (.A ( n1409 ) , .B ( n1408 ) , .Y ( n1410 ));
INVX2 U1409  (.A ( n1508 ) , .Y ( n1509 ));
CLKXOR2X4 U1410  (.A ( n1811 ) , .B ( n1804 ) , .Y ( n1854 ));
XOR2X1 U1411  (.A ( n1838 ) , .B ( n1839 ) , .Y ( n1829 ));
NAND2X4 U1412  (.A ( n1556 ) , .B ( \intadd_7/SUM[2] ) , .Y ( n1699 ));
NAND2X4 U1413  (.A ( n1373 ) , .B ( n1372 ) , .Y ( n1382 ));
NAND2X4 U1414  (.A ( n1517 ) , .B ( n1558 ) , .Y ( n1568 ));
INVX2 U1415  (.A ( n1371 ) , .Y ( n1372 ));
NAND2X2 U1416  (.A ( n1790 ) , .B ( n1788 ) , .Y ( n1805 ));
XOR2X1 U1417  (.A ( n1813 ) , .B ( n1797 ) , .Y ( n1798 ));
NAND2BX8 U1418  (.AN ( n1726 ) , .B ( n1725 ) , .Y ( n1767 ));
INVX2 U1419  (.A ( n1765 ) , .Y ( n1766 ));
NAND2X2 U1420  (.A ( n1357 ) , .B ( n1338 ) , .Y ( n1194 ));
NAND2X2 U1421  (.A ( n1283 ) , .B ( n1453 ) , .Y ( n1299 ));
NAND2X2 U1422  (.A ( n1794 ) , .B ( a[6] ) , .Y ( n1795 ));
INVX2 U1423  (.A ( n1455 ) , .Y ( n1283 ));
INVXL U1424  (.A ( n1647 ) , .Y ( n1601 ));
XOR2XL U1425  (.A ( n1648 ) , .B ( n1649 ) , .Y ( n1602 ));
OAI21X2 U1426  (.A0 ( n1625 ) , .A1 ( n1624 ) , .B0 ( n1623 ) , .Y ( n1627 ));
XOR2X2 U1427  (.A ( n1295 ) , .B ( n1294 ) , .Y ( n1354 ));
INVX4 U1428  (.A ( n2742 ) , .Y ( n2305 ));
NAND2X4 U1429  (.A ( n1181 ) , .B ( n1180 ) , .Y ( n1300 ));
AOI21X2 U1430  (.A0 ( n2754 ) , .A1 ( n1280 ) , .B0 ( \intadd_7/A[0] ) , .Y ( n1281 ));
OAI21X2 U1431  (.A0 ( n1209 ) , .A1 ( n1208 ) , .B0 ( n1212 ) , .Y ( n1232 ));
INVX2 U1432  (.A ( n1741 ) , .Y ( n1742 ));
NAND2X2 U1433  (.A ( n1613 ) , .B ( n1612 ) , .Y ( n2752 ));
XOR2X2 U1434  (.A ( n1157 ) , .B ( n1156 ) , .Y ( n1158 ));
NAND2X2 U1435  (.A ( n1348 ) , .B ( n1347 ) , .Y ( n1349 ));
INVX1 U1436  (.A ( n1219 ) , .Y ( n1204 ));
NAND2X2 U1437  (.A ( n1716 ) , .B ( n2733 ) , .Y ( n1656 ));
AND2XL U1438  (.A ( n2029 ) , .B ( n2028 ) , .Y ( n2032 ));
XOR2XL U1439  (.A ( n2120 ) , .B ( n2119 ) , .Y ( n2121 ));
NAND2X2 U1440  (.A ( n1707 ) , .B ( n1121 ) , .Y ( n1187 ));
NAND2X2 U1441  (.A ( n1750 ) , .B ( n1834 ) , .Y ( n1782 ));
XOR2XL U1442  (.A ( n1234 ) , .B ( n1233 ) , .Y ( n1236 ));
INVX1 U1443  (.A ( n2754 ) , .Y ( n2757 ));
INVXL U1444  (.A ( n1424 ) , .Y ( n1425 ));
INVX2 U1445  (.A ( n1839 ) , .Y ( n1840 ));
OAI2BB1XL U1446  (.A0N ( n1049 ) , .A1N ( n1866 ) , .B0 ( n1865 ) , .Y ( n1868 ));
NAND2BXL U1447  (.AN ( n1865 ) , .B ( n1049 ) , .Y ( n1848 ));
NAND2X1 U1448  (.A ( n2008 ) , .B ( n2009 ) , .Y ( n2012 ));
INVX2 U1449  (.A ( n1353 ) , .Y ( n1288 ));
NAND2X1 U1450  (.A ( n2734 ) , .B ( n2702 ) , .Y ( n1611 ));
INVX2 U1451  (.A ( n1491 ) , .Y ( n1495 ));
NAND2XL U1452  (.A ( n1976 ) , .B ( n1972 ) , .Y ( n1967 ));
MXI2X2 U1453  (.A ( n1251 ) , .B ( n1250 ) , .S0 ( n1403 ) , .Y ( n1252 ));
INVX2 U1454  (.A ( n1846 ) , .Y ( n1866 ));
INVXL U1455  (.A ( n1231 ) , .Y ( n1210 ));
NAND2X4 U1456  (.A ( n1063 ) , .B ( n1877 ) , .Y ( n1091 ));
NAND2X2 U1457  (.A ( n1490 ) , .B ( n2731 ) , .Y ( n1268 ));
NAND2X2 U1458  (.A ( n1974 ) , .B ( \intadd_4/n1  ) , .Y ( n1083 ));
NAND2X2 U1459  (.A ( n2699 ) , .B ( n2702 ) , .Y ( n2700 ));
NAND2XL U1460  (.A ( n1920 ) , .B ( n1956 ) , .Y ( n1941 ));
NAND2X2 U1461  (.A ( n1492 ) , .B ( n1820 ) , .Y ( n1541 ));
NAND2X4 U1462  (.A ( n1820 ) , .B ( n1818 ) , .Y ( n1799 ));
INVX2 U1463  (.A ( n1062 ) , .Y ( n1060 ));
NAND2X2 U1464  (.A ( n2702 ) , .B ( n2750 ) , .Y ( n1186 ));
NOR2X4 U1465  (.A ( n1049 ) , .B ( n1403 ) , .Y ( n1412 ));
INVX12 U1466  (.A ( n1088 ) , .Y ( n1093 ));
NAND4BXL U1467  (.AN ( b[10] ) , .B ( n1875 ) , .C ( n1874 ) , .D ( n2761 ) , .Y ( n1876 ));
INVX4 U1468  (.A ( b[3] ) , .Y ( n1109 ));
INVX2 U1469  (.A ( c[14] ) , .Y ( n1984 ));
AND2XL U1470  (.A ( a[10] ) , .B ( b[10] ) , .Y ( \intadd_4/CI  ));
INVXL U1471  (.A ( c[15] ) , .Y ( n2291 ));
OAI21X4 U1472  (.A0 ( n2501 ) , .A1 ( n2651 ) , .B0 ( n1054 ) , .Y ( n2502 ));
XOR2X2 U1473  (.A ( n2602 ) , .B ( n2601 ) , .Y ( n2604 ));
INVX4 U1474  (.A ( n2603 ) , .Y ( n2514 ));
CLKNAND2X12 U1475  (.A ( n2556 ) , .B ( n2474 ) , .Y ( n2671 ));
XOR2X2 U1476  (.A ( n2642 ) , .B ( n2600 ) , .Y ( n2602 ));
AOI211X2 U1477  (.A0 ( n2626 ) , .A1 ( n2625 ) , .B0 ( n2624 ) , .C0 ( n2742 ) , .Y ( n2630 ));
INVX2 U1478  (.A ( n2686 ) , .Y ( n2500 ));
NAND2X4 U1479  (.A ( n2623 ) , .B ( n2543 ) , .Y ( n2512 ));
NOR4X2 U1480  (.A ( n2726 ) , .B ( n2725 ) , .C ( n2724 ) , .D ( n2655 ) , .Y ( n2607 ));
OAI22X2 U1481  (.A0 ( n2668 ) , .A1 ( n2544 ) , .B0 ( n2628 ) , .B1 ( n2543 ) , .Y ( n2545 ));
OR2X2 U1482  (.A ( n2650 ) , .B ( n2694 ) , .Y ( n1054 ));
INVX4 U1483  (.A ( n2678 ) , .Y ( n2666 ));
NOR2X2 U1484  (.A ( n2628 ) , .B ( n2598 ) , .Y ( n2724 ));
AND3X6 U1485  (.A ( n2454 ) , .B ( n2591 ) , .C ( n2588 ) , .Y ( n2508 ));
INVX2 U1486  (.A ( n2588 ) , .Y ( n2631 ));
NOR2X2 U1487  (.A ( n2542 ) , .B ( n2556 ) , .Y ( n2546 ));
XNOR2X1 U1488  (.A ( n2563 ) , .B ( n2567 ) , .Y ( n2565 ));
AOI21X4 U1489  (.A0 ( n2519 ) , .A1 ( n2548 ) , .B0 ( n2562 ) , .Y ( n2520 ));
NAND3X4 U1490  (.A ( n2465 ) , .B ( n2467 ) , .C ( n2464 ) , .Y ( n2472 ));
XOR2X4 U1491  (.A ( n2409 ) , .B ( n2408 ) , .Y ( n2677 ));
INVX4 U1492  (.A ( n2694 ) , .Y ( n2584 ));
XOR2X4 U1493  (.A ( n2400 ) , .B ( n2433 ) , .Y ( n2694 ));
NAND3X6 U1494  (.A ( n2399 ) , .B ( n2398 ) , .C ( n2406 ) , .Y ( n2433 ));
NAND2BX4 U1495  (.AN ( n2304 ) , .B ( n2302 ) , .Y ( n2434 ));
INVX2 U1496  (.A ( n2422 ) , .Y ( n2405 ));
NAND2X4 U1497  (.A ( n2299 ) , .B ( n2298 ) , .Y ( n2304 ));
INVX4 U1498  (.A ( n2385 ) , .Y ( n2388 ));
NAND2X4 U1499  (.A ( n2385 ) , .B ( n2386 ) , .Y ( n2423 ));
NAND2X4 U1500  (.A ( n2429 ) , .B ( n2456 ) , .Y ( n2403 ));
INVX2 U1501  (.A ( n2455 ) , .Y ( n2427 ));
NAND2X4 U1502  (.A ( n2492 ) , .B ( n2493 ) , .Y ( n2354 ));
NAND3X4 U1503  (.A ( n2370 ) , .B ( n2305 ) , .C ( n2369 ) , .Y ( n2394 ));
NAND2X4 U1504  (.A ( n2328 ) , .B ( n2358 ) , .Y ( n2331 ));
NAND2X4 U1505  (.A ( n2363 ) , .B ( n2364 ) , .Y ( n2455 ));
NAND3X4 U1506  (.A ( n2312 ) , .B ( n2311 ) , .C ( n2310 ) , .Y ( n2363 ));
NAND2X4 U1507  (.A ( n2478 ) , .B ( n2477 ) , .Y ( n2658 ));
MXI2X2 U1508  (.A ( n2334 ) , .B ( n2338 ) , .S0 ( n2333 ) , .Y ( n2336 ));
INVX2 U1509  (.A ( n2389 ) , .Y ( n2392 ));
AND2X6 U1510  (.A ( n2257 ) , .B ( n2256 ) , .Y ( n2340 ));
AOI21X4 U1511  (.A0 ( n2202 ) , .A1 ( n2283 ) , .B0 ( n2201 ) , .Y ( n2206 ));
INVX2 U1512  (.A ( n2442 ) , .Y ( n2443 ));
INVX2 U1513  (.A ( n2308 ) , .Y ( n2306 ));
NAND3X4 U1514  (.A ( n2234 ) , .B ( n2286 ) , .C ( n2235 ) , .Y ( n2230 ));
NAND2X4 U1515  (.A ( n2273 ) , .B ( n2411 ) , .Y ( n2324 ));
NAND3X4 U1516  (.A ( n2410 ) , .B ( n2235 ) , .C ( n2234 ) , .Y ( n2257 ));
NAND2X6 U1517  (.A ( n2411 ) , .B ( n2286 ) , .Y ( n2297 ));
NOR2X6 U1518  (.A ( n2259 ) , .B ( n2266 ) , .Y ( n2410 ));
NAND2BX2 U1519  (.AN ( n2269 ) , .B ( n2265 ) , .Y ( n2261 ));
NAND2X2 U1520  (.A ( n2278 ) , .B ( n2274 ) , .Y ( n2262 ));
NAND2X6 U1521  (.A ( n2221 ) , .B ( n2275 ) , .Y ( n2259 ));
NAND2X6 U1522  (.A ( n2275 ) , .B ( n2193 ) , .Y ( n2439 ));
NAND2X4 U1523  (.A ( n2179 ) , .B ( n2178 ) , .Y ( n2196 ));
AOI21X6 U1524  (.A0 ( n2195 ) , .A1 ( n2199 ) , .B0 ( n2186 ) , .Y ( n2252 ));
NAND2X4 U1525  (.A ( n2203 ) , .B ( n2280 ) , .Y ( n2247 ));
MXI2X2 U1526  (.A ( n2279 ) , .B ( n2277 ) , .S0 ( n2280 ) , .Y ( n2229 ));
INVX2 U1527  (.A ( n2266 ) , .Y ( n2267 ));
INVX2 U1528  (.A ( n2302 ) , .Y ( n2303 ));
INVX2 U1529  (.A ( n2268 ) , .Y ( n2260 ));
MXI2X1 U1530  (.A ( n2248 ) , .B ( n2242 ) , .S0 ( n2277 ) , .Y ( n2209 ));
MXI2X1 U1531  (.A ( c[6] ) , .B ( n2382 ) , .S0 ( n2621 ) , .Y ( n2386 ));
INVX1 U1532  (.A ( n2236 ) , .Y ( n2240 ));
INVX2 U1533  (.A ( n2232 ) , .Y ( n2233 ));
MXI2XL U1534  (.A ( n2483 ) , .B ( n2346 ) , .S0 ( n2218 ) , .Y ( n2220 ));
MXI2X1 U1535  (.A ( c[1] ) , .B ( n2348 ) , .S0 ( n2218 ) , .Y ( n2236 ));
MXI2X2 U1536  (.A ( c[7] ) , .B ( n2372 ) , .S0 ( n2218 ) , .Y ( n2246 ));
MXI2X4 U1537  (.A ( c[13] ) , .B ( n2527 ) , .S0 ( n2189 ) , .Y ( n2184 ));
NOR2X2 U1538  (.A ( n2553 ) , .B ( n2551 ) , .Y ( n2610 ));
NOR2X2 U1539  (.A ( n2525 ) , .B ( n2524 ) , .Y ( n2551 ));
INVX2 U1540  (.A ( n2463 ) , .Y ( n2468 ));
INVX2 U1541  (.A ( n2151 ) , .Y ( n2153 ));
NOR2X2 U1542  (.A ( n2528 ) , .B ( n2556 ) , .Y ( n2530 ));
INVX1 U1543  (.A ( n2567 ) , .Y ( n2740 ));
NOR2X2 U1544  (.A ( n2555 ) , .B ( n2556 ) , .Y ( n2558 ));
NAND3X4 U1545  (.A ( n2135 ) , .B ( n2540 ) , .C ( n2548 ) , .Y ( n2140 ));
NAND2X4 U1546  (.A ( n2527 ) , .B ( n2537 ) , .Y ( n2139 ));
NOR2X2 U1547  (.A ( n2445 ) , .B ( n2556 ) , .Y ( n2463 ));
NAND2X4 U1548  (.A ( n1971 ) , .B ( n1970 ) , .Y ( n1983 ));
NAND2X4 U1549  (.A ( n1943 ) , .B ( n1942 ) , .Y ( n1944 ));
AND3X6 U1550  (.A ( n2126 ) , .B ( n2125 ) , .C ( n2124 ) , .Y ( n2187 ));
NAND2BX4 U1551  (.AN ( n2211 ) , .B ( n1919 ) , .Y ( n1916 ));
AOI21X4 U1552  (.A0 ( n2116 ) , .A1 ( n2115 ) , .B0 ( n2114 ) , .Y ( n2122 ));
NAND2X4 U1553  (.A ( n2084 ) , .B ( n2083 ) , .Y ( n2110 ));
AND2X4 U1554  (.A ( n1935 ) , .B ( n2076 ) , .Y ( n1977 ));
NAND2X2 U1555  (.A ( n2016 ) , .B ( n1936 ) , .Y ( n1935 ));
AND2X4 U1556  (.A ( n1773 ) , .B ( n1772 ) , .Y ( n1891 ));
INVX1 U1557  (.A ( n1994 ) , .Y ( n1995 ));
INVX4 U1558  (.A ( n1668 ) , .Y ( n1664 ));
NAND3X6 U1559  (.A ( n1740 ) , .B ( n1739 ) , .C ( n1738 ) , .Y ( n1755 ));
INVX2 U1560  (.A ( n1927 ) , .Y ( n1930 ));
INVX2 U1561  (.A ( n2108 ) , .Y ( n1911 ));
NAND2X4 U1562  (.A ( n1734 ) , .B ( n1733 ) , .Y ( n1735 ));
INVX2 U1563  (.A ( n2103 ) , .Y ( n2107 ));
AND2X4 U1564  (.A ( n1728 ) , .B ( n1732 ) , .Y ( n1737 ));
INVX4 U1565  (.A ( n1499 ) , .Y ( n1484 ));
INVX2 U1566  (.A ( n1444 ) , .Y ( n1447 ));
NAND2X2 U1567  (.A ( n1677 ) , .B ( n1692 ) , .Y ( n1691 ));
AND3X2 U1568  (.A ( n2097 ) , .B ( c[8] ) , .C ( n2095 ) , .Y ( n2089 ));
OAI21X6 U1569  (.A0 ( n1573 ) , .A1 ( n1572 ) , .B0 ( n1693 ) , .Y ( n1588 ));
AND2X4 U1570  (.A ( n1385 ) , .B ( n1384 ) , .Y ( n1407 ));
INVX2 U1571  (.A ( n1774 ) , .Y ( n1775 ));
NAND2X2 U1572  (.A ( n1808 ) , .B ( n1807 ) , .Y ( n1809 ));
NAND2X2 U1573  (.A ( n1699 ) , .B ( n1569 ) , .Y ( n1559 ));
XOR2X1 U1574  (.A ( n1803 ) , .B ( n1810 ) , .Y ( n1804 ));
NAND2X6 U1575  (.A ( n1395 ) , .B ( n1394 ) , .Y ( n1405 ));
AND2X2 U1576  (.A ( n1221 ) , .B ( n1224 ) , .Y ( n1052 ));
INVX2 U1577  (.A ( n1807 ) , .Y ( n1803 ));
INVX2 U1578  (.A ( n1813 ) , .Y ( n1814 ));
NAND3X2 U1579  (.A ( n1696 ) , .B ( n1695 ) , .C ( n1694 ) , .Y ( n1697 ));
XOR2X2 U1580  (.A ( n1743 ) , .B ( n1741 ) , .Y ( n1694 ));
NAND2X4 U1581  (.A ( n1724 ) , .B ( n1723 ) , .Y ( n1726 ));
NAND2X2 U1582  (.A ( n1515 ) , .B ( n1513 ) , .Y ( n1462 ));
AOI21X1 U1583  (.A0 ( n1344 ) , .A1 ( n1343 ) , .B0 ( n1342 ) , .Y ( n1345 ));
OAI21X4 U1584  (.A0 ( n1684 ) , .A1 ( n1683 ) , .B0 ( n1682 ) , .Y ( n1743 ));
XOR2X2 U1585  (.A ( n1199 ) , .B ( n1198 ) , .Y ( n1200 ));
CLKXOR2X4 U1586  (.A ( n1794 ) , .B ( n1764 ) , .Y ( n1765 ));
INVX2 U1587  (.A ( n1366 ) , .Y ( n1298 ));
INVX1 U1588  (.A ( n2051 ) , .Y ( n1244 ));
OAI21X2 U1589  (.A0 ( n1681 ) , .A1 ( n1680 ) , .B0 ( n1679 ) , .Y ( n1682 ));
INVXL U1590  (.A ( n1725 ) , .Y ( n1727 ));
ADDFX2 U1591  (.A ( \intadd_7/A[2] ) , .B ( \intadd_7/B[2] ) , .CI ( \intadd_7/n2  ) , .CO ( \intadd_7/n1  ) , .S ( \intadd_7/SUM[2] ));
INVX2 U1592  (.A ( n1587 ) , .Y ( n1585 ));
OAI21X2 U1593  (.A0 ( n1649 ) , .A1 ( n1648 ) , .B0 ( n1647 ) , .Y ( n1650 ));
INVXL U1594  (.A ( n1721 ) , .Y ( n1661 ));
NAND2X4 U1595  (.A ( n1627 ) , .B ( n1626 ) , .Y ( n1681 ));
INVX2 U1596  (.A ( n2037 ) , .Y ( n1243 ));
NAND2X2 U1597  (.A ( n1302 ) , .B ( n1300 ) , .Y ( n1192 ));
INVX2 U1598  (.A ( n1198 ) , .Y ( n1167 ));
NAND2BX2 U1599  (.AN ( n1832 ) , .B ( n1831 ) , .Y ( n1833 ));
INVX2 U1600  (.A ( n1532 ) , .Y ( n1533 ));
NOR2X2 U1601  (.A ( n1354 ) , .B ( n1353 ) , .Y ( n1355 ));
INVX4 U1602  (.A ( n2305 ) , .Y ( n2550 ));
INVX2 U1603  (.A ( n1812 ) , .Y ( n1815 ));
OAI21X4 U1604  (.A0 ( n1597 ) , .A1 ( n1596 ) , .B0 ( n1595 ) , .Y ( n1654 ));
INVX2 U1605  (.A ( n2710 ) , .Y ( n2703 ));
NAND2X4 U1606  (.A ( n1546 ) , .B ( n1545 ) , .Y ( n1649 ));
NAND2BX2 U1607  (.AN ( n1812 ) , .B ( n2702 ) , .Y ( n1797 ));
XOR2X2 U1608  (.A ( n1159 ) , .B ( n1158 ) , .Y ( n1213 ));
NAND2X4 U1609  (.A ( n1154 ) , .B ( n1153 ) , .Y ( n1181 ));
AOI21X4 U1610  (.A0 ( n1256 ) , .A1 ( n1255 ) , .B0 ( n1254 ) , .Y ( n1294 ));
NOR2X4 U1611  (.A ( n2705 ) , .B ( n2704 ) , .Y ( n2710 ));
CLKXOR2X2 U1612  (.A ( n1631 ) , .B ( n1583 ) , .Y ( n1620 ));
INVX2 U1613  (.A ( n1714 ) , .Y ( n1718 ));
NAND2BX2 U1614  (.AN ( n1715 ) , .B ( n1706 ) , .Y ( n1658 ));
NAND2X2 U1615  (.A ( n1256 ) , .B ( n1253 ) , .Y ( n1105 ));
OAI21X2 U1616  (.A0 ( n1540 ) , .A1 ( n1539 ) , .B0 ( n1538 ) , .Y ( n1592 ));
NOR2X2 U1617  (.A ( n2708 ) , .B ( n2707 ) , .Y ( n2709 ));
OAI21X4 U1618  (.A0 ( n1142 ) , .A1 ( n1161 ) , .B0 ( n1141 ) , .Y ( n1144 ));
NOR2X2 U1619  (.A ( n1280 ) , .B ( n2754 ) , .Y ( \intadd_7/A[0] ));
CLKXOR2X2 U1620  (.A ( n1579 ) , .B ( n1529 ) , .Y ( n1530 ));
INVX2 U1621  (.A ( n1480 ) , .Y ( n1478 ));
INVX4 U1622  (.A ( n1162 ) , .Y ( n1141 ));
INVX2 U1623  (.A ( n2755 ) , .Y ( n1616 ));
AND2X4 U1624  (.A ( n1319 ) , .B ( n1178 ) , .Y ( n1179 ));
NAND2BX2 U1625  (.AN ( n1712 ) , .B ( n2702 ) , .Y ( n1713 ));
INVX2 U1626  (.A ( n1862 ) , .Y ( n1863 ));
NOR2X2 U1627  (.A ( n2698 ) , .B ( n1091 ) , .Y ( n2701 ));
NAND2X2 U1628  (.A ( n1748 ) , .B ( n1749 ) , .Y ( n1746 ));
NOR2X2 U1629  (.A ( n2756 ) , .B ( n2732 ) , .Y ( n1614 ));
NAND2BX2 U1630  (.AN ( n1652 ) , .B ( n1653 ) , .Y ( n1600 ));
OAI22X1 U1631  (.A0 ( n1177 ) , .A1 ( n1474 ) , .B0 ( n1176 ) , .B1 ( n1175 ) , .Y ( n1178 ));
NOR2X2 U1632  (.A ( n1255 ) , .B ( n1203 ) , .Y ( n1219 ));
OR2X2 U1633  (.A ( error ) , .B ( n2289 ) , .Y ( n1057 ));
NAND2BX2 U1634  (.AN ( n2289 ) , .B ( n2288 ) , .Y ( n2619 ));
INVX1 U1635  (.A ( n2012 ) , .Y ( n1987 ));
NOR2X2 U1636  (.A ( n1706 ) , .B ( n1800 ) , .Y ( n1546 ));
INVX2 U1637  (.A ( n1156 ) , .Y ( n1147 ));
NOR2X2 U1638  (.A ( n1830 ) , .B ( n1786 ) , .Y ( n1787 ));
NOR2X2 U1639  (.A ( n1272 ) , .B ( n1257 ) , .Y ( n1258 ));
BUFX10 U1640  (.A ( n1068 ) , .Y ( n2733 ));
NAND2BX2 U1641  (.AN ( n1685 ) , .B ( n1632 ) , .Y ( n1634 ));
OAI21X3 U1642  (.A0 ( n1172 ) , .A1 ( n1170 ) , .B0 ( n1114 ) , .Y ( n1115 ));
AOI21X4 U1643  (.A0 ( n1135 ) , .A1 ( n1133 ) , .B0 ( n1124 ) , .Y ( n1156 ));
XOR2X2 U1644  (.A ( n1076 ) , .B ( n1075 ) , .Y ( n1077 ));
XOR2X2 U1645  (.A ( n1067 ) , .B ( n1759 ) , .Y ( n1068 ));
NAND2X4 U1646  (.A ( n1252 ) , .B ( n1472 ) , .Y ( n1522 ));
NAND2X4 U1647  (.A ( n1882 ) , .B ( n1093 ) , .Y ( n1076 ));
NAND2BX2 U1648  (.AN ( n1091 ) , .B ( n2702 ) , .Y ( n2707 ));
INVXL U1649  (.A ( n1091 ) , .Y ( n1289 ));
AND2X1 U1650  (.A ( n2004 ) , .B ( n2020 ) , .Y ( n2009 ));
INVX4 U1651  (.A ( n1148 ) , .Y ( n1170 ));
AOI21X1 U1652  (.A0 ( n2118 ) , .A1 ( n1820 ) , .B0 ( n1819 ) , .Y ( n1821 ));
NOR2X2 U1653  (.A ( n1802 ) , .B ( n1403 ) , .Y ( n1433 ));
AOI21X4 U1654  (.A0 ( n1060 ) , .A1 ( n1059 ) , .B0 ( n1058 ) , .Y ( n1063 ));
INVX4 U1655  (.A ( n1799 ) , .Y ( n1657 ));
NAND2X2 U1656  (.A ( n2731 ) , .B ( n2748 ) , .Y ( n1101 ));
OR2X2 U1657  (.A ( n1492 ) , .B ( n2748 ) , .Y ( n1490 ));
INVX2 U1658  (.A ( n1593 ) , .Y ( n1597 ));
NOR2X2 U1659  (.A ( n1918 ) , .B ( n1957 ) , .Y ( n1942 ));
MXI2X2 U1660  (.A ( n1094 ) , .B ( n1093 ) , .S0 ( n2760 ) , .Y ( n1096 ));
INVX6 U1661  (.A ( n1092 ) , .Y ( n1065 ));
AND2X2 U1662  (.A ( a[1] ) , .B ( n2556 ) , .Y ( n1536 ));
AND2X6 U1663  (.A ( n2556 ) , .B ( b[9] ) , .Y ( n1818 ));
NAND2BX2 U1664  (.AN ( n2556 ) , .B ( c[10] ) , .Y ( n2461 ));
NOR2X6 U1665  (.A ( n1069 ) , .B ( b[4] ) , .Y ( n1062 ));
NOR2X4 U1666  (.A ( n1088 ) , .B ( n1430 ) , .Y ( n1089 ));
NAND2X4 U1667  (.A ( n1064 ) , .B ( n1085 ) , .Y ( n1092 ));
NOR2X6 U1668  (.A ( n1112 ) , .B ( b[2] ) , .Y ( n1106 ));
INVX12 U1669  (.A ( n2643 ) , .Y ( n2293 ));
NAND4BX2 U1670  (.AN ( a[10] ) , .B ( n1880 ) , .C ( n1879 ) , .D ( n1878 ) , .Y ( n1881 ));
AND2XL U1671  (.A ( c[11] ) , .B ( c[10] ) , .Y ( n2158 ));
BUFX8 U1672  (.A ( n2749 ) , .Y ( n1048 ));
OAI211X2 U1673  (.A0 ( n2738 ) , .A1 ( n2576 ) , .B0 ( n2575 ) , .C0 ( n2574 ) , .Y ( n997 ));
NAND2BX2 U1674  (.AN ( n2736 ) , .B ( n2518 ) , .Y ( n2534 ));
MXI2X1 U1675  (.A ( n2715 ) , .B ( n2503 ) , .S0 ( n2655 ) , .Y ( n1004 ));
MXI2X1 U1676  (.A ( n2711 ) , .B ( n2664 ) , .S0 ( n2655 ) , .Y ( n1008 ));
MXI2X1 U1677  (.A ( n2717 ) , .B ( n2656 ) , .S0 ( n2655 ) , .Y ( n1006 ));
MXI2X2 U1678  (.A ( n2645 ) , .B ( n2644 ) , .S0 ( n2643 ) , .Y ( n2716 ));
MXI2X1 U1679  (.A ( n2713 ) , .B ( n2548 ) , .S0 ( n2655 ) , .Y ( n1000 ));
NOR4X4 U1680  (.A ( n2571 ) , .B ( n2570 ) , .C ( n2549 ) , .D ( n2550 ) , .Y ( n2518 ));
INVX4 U1681  (.A ( n2671 ) , .Y ( n2695 ));
XOR2X4 U1682  (.A ( n2604 ) , .B ( n2603 ) , .Y ( n2722 ));
MXI2X1 U1683  (.A ( n2714 ) , .B ( n2632 ) , .S0 ( n2655 ) , .Y ( n1001 ));
AOI22X2 U1684  (.A0 ( n2589 ) , .A1 ( n2690 ) , .B0 ( n2689 ) , .B1 ( n2631 ) , .Y ( n2590 ));
AOI21X4 U1685  (.A0 ( n2500 ) , .A1 ( n2670 ) , .B0 ( n2499 ) , .Y ( n2501 ));
AOI22X2 U1686  (.A0 ( n2570 ) , .A1 ( n2517 ) , .B0 ( n2507 ) , .B1 ( n2506 ) , .Y ( n2536 ));
OAI22X2 U1687  (.A0 ( n2745 ) , .A1 ( n2566 ) , .B0 ( c[14] ) , .B1 ( n2749 ) , .Y ( n2575 ));
OAI21X1 U1688  (.A0 ( n2633 ) , .A1 ( n2658 ) , .B0 ( n2578 ) , .Y ( n2579 ));
NAND3BX2 U1689  (.AN ( n2587 ) , .B ( n2586 ) , .C ( n2585 ) , .Y ( n2589 ));
OAI22X2 U1690  (.A0 ( n2620 ) , .A1 ( n2556 ) , .B0 ( n2218 ) , .B1 ( n2619 ) , .Y ( n2728 ));
XOR2X1 U1691  (.A ( n2618 ) , .B ( n2651 ) , .Y ( n2620 ));
NOR2X6 U1692  (.A ( n2623 ) , .B ( n2543 ) , .Y ( n2511 ));
AOI2BB2X1 U1693  (.B0 ( n2666 ) , .B1 ( n2584 ) , .A0N ( n2686 ) , .A1N ( n2679 ) , .Y ( n2585 ));
XNOR2X1 U1694  (.A ( n2533 ) , .B ( n2532 ) , .Y ( n1050 ));
AOI21X1 U1695  (.A0 ( n2617 ) , .A1 ( n2593 ) , .B0 ( n2526 ) , .Y ( n2533 ));
BUFX10 U1696  (.A ( n2460 ) , .Y ( n2674 ));
OAI21X1 U1697  (.A0 ( n2668 ) , .A1 ( n2561 ) , .B0 ( n2568 ) , .Y ( n2506 ));
MXI2X1 U1698  (.A ( n2668 ) , .B ( n2628 ) , .S0 ( n2627 ) , .Y ( n2629 ));
OAI22X1 U1699  (.A0 ( n2680 ) , .A1 ( n2658 ) , .B0 ( n2647 ) , .B1 ( n2678 ) , .Y ( n2648 ));
XOR2X1 U1700  (.A ( n2562 ) , .B ( n2541 ) , .Y ( n2542 ));
NAND2X4 U1701  (.A ( n2438 ) , .B ( n2437 ) , .Y ( n2450 ));
AND3X4 U1702  (.A ( n2432 ) , .B ( n2673 ) , .C ( n2654 ) , .Y ( n2451 ));
XOR2X2 U1703  (.A ( n2434 ) , .B ( n2452 ) , .Y ( n2432 ));
INVX4 U1704  (.A ( n2466 ) , .Y ( n2437 ));
NAND2BX4 U1705  (.AN ( n2421 ) , .B ( n2420 ) , .Y ( n2465 ));
NAND2X4 U1706  (.A ( n2304 ) , .B ( n2303 ) , .Y ( n2435 ));
NAND2X4 U1707  (.A ( n2444 ) , .B ( n2414 ) , .Y ( n2417 ));
NAND2X4 U1708  (.A ( n2388 ) , .B ( n2387 ) , .Y ( n2422 ));
OAI21X6 U1709  (.A0 ( n2362 ) , .A1 ( n2378 ) , .B0 ( n2361 ) , .Y ( n2429 ));
NAND2BX4 U1710  (.AN ( n2378 ) , .B ( n2377 ) , .Y ( n2379 ));
INVX4 U1711  (.A ( n2356 ) , .Y ( n2323 ));
NAND2X4 U1712  (.A ( n2481 ) , .B ( n2479 ) , .Y ( n2350 ));
NAND2X4 U1713  (.A ( n2336 ) , .B ( n2335 ) , .Y ( n2353 ));
AOI21X6 U1714  (.A0 ( n2320 ) , .A1 ( n2319 ) , .B0 ( n2318 ) , .Y ( n2356 ));
INVX1 U1715  (.A ( n2333 ) , .Y ( n2316 ));
INVX4 U1716  (.A ( n2324 ) , .Y ( n2327 ));
NAND3X4 U1717  (.A ( n2263 ) , .B ( n2262 ) , .C ( n2261 ) , .Y ( n2264 ));
NAND3X4 U1718  (.A ( n2228 ) , .B ( n2227 ) , .C ( n2226 ) , .Y ( n2231 ));
NAND2X4 U1719  (.A ( n2196 ) , .B ( n2195 ) , .Y ( n2198 ));
INVX12 U1720  (.A ( n2203 ) , .Y ( n2275 ));
NOR2X4 U1721  (.A ( n2280 ) , .B ( n2277 ) , .Y ( n2193 ));
NAND2X6 U1722  (.A ( n2174 ) , .B ( n2568 ) , .Y ( n2195 ));
NAND2BX4 U1723  (.AN ( n2177 ) , .B ( n2179 ) , .Y ( n2164 ));
OAI21X1 U1724  (.A0 ( n2729 ) , .A1 ( n2655 ) , .B0 ( c[15] ) , .Y ( n2622 ));
NAND2X4 U1725  (.A ( n2183 ) , .B ( n2173 ) , .Y ( n2174 ));
AOI21X6 U1726  (.A0 ( n2156 ) , .A1 ( n2172 ) , .B0 ( n2601 ) , .Y ( n2177 ));
MXI2X1 U1727  (.A ( c[7] ) , .B ( n2372 ) , .S0 ( n2621 ) , .Y ( n2395 ));
MXI2X1 U1728  (.A ( n2243 ) , .B ( n2242 ) , .S0 ( n2241 ) , .Y ( n2258 ));
INVX1 U1729  (.A ( n2621 ) , .Y ( n2729 ));
MXI2X1 U1730  (.A ( c[0] ) , .B ( n2347 ) , .S0 ( n2621 ) , .Y ( n2476 ));
INVX1 U1731  (.A ( n2601 ) , .Y ( n2598 ));
AND2X4 U1732  (.A ( n2504 ) , .B ( n2163 ) , .Y ( n2165 ));
OAI21X6 U1733  (.A0 ( n2134 ) , .A1 ( n2133 ) , .B0 ( n2132 ) , .Y ( n2145 ));
OAI21X1 U1734  (.A0 ( n2553 ) , .A1 ( n2592 ) , .B0 ( n2552 ) , .Y ( n2614 ));
INVX1 U1735  (.A ( n2551 ) , .Y ( n2593 ));
NOR2X4 U1736  (.A ( n1986 ) , .B ( n1985 ) , .Y ( n2146 ));
NAND2X1 U1737  (.A ( n2530 ) , .B ( n2529 ) , .Y ( n2552 ));
AND2X1 U1738  (.A ( n2740 ) , .B ( n2599 ) , .Y ( n2572 ));
OAI21X2 U1739  (.A0 ( n2527 ) , .A1 ( n2537 ) , .B0 ( n2182 ) , .Y ( n2143 ));
NAND4X4 U1740  (.A ( n2101 ) , .B ( n2127 ) , .C ( n2646 ) , .D ( n2382 ) , .Y ( n2130 ));
NAND2BX4 U1741  (.AN ( n2554 ) , .B ( n1051 ) , .Y ( n2182 ));
NAND2X8 U1742  (.A ( n1969 ) , .B ( n1968 ) , .Y ( n2527 ));
INVXL U1743  (.A ( n2329 ) , .Y ( n2330 ));
INVXL U1744  (.A ( n2313 ) , .Y ( n2314 ));
NAND3X6 U1745  (.A ( n2032 ) , .B ( n2031 ) , .C ( n2030 ) , .Y ( n2337 ));
AND3X1 U1746  (.A ( n2217 ) , .B ( n2216 ) , .C ( n2215 ) , .Y ( n2346 ));
NAND3X6 U1747  (.A ( n2061 ) , .B ( n2060 ) , .C ( n2059 ) , .Y ( n2329 ));
NAND2BX4 U1748  (.AN ( n2214 ) , .B ( n2102 ) , .Y ( n2098 ));
XOR2X4 U1749  (.A ( n1902 ) , .B ( n1901 ) , .Y ( n2079 ));
AOI21X6 U1750  (.A0 ( n2116 ) , .A1 ( n2085 ) , .B0 ( n2110 ) , .Y ( n2088 ));
AOI21X6 U1751  (.A0 ( n2116 ) , .A1 ( n2080 ) , .B0 ( n1900 ) , .Y ( n1902 ));
NAND3X6 U1752  (.A ( n1893 ) , .B ( n1892 ) , .C ( n2041 ) , .Y ( n2057 ));
NAND3X4 U1753  (.A ( n1778 ) , .B ( n1777 ) , .C ( n2056 ) , .Y ( n1851 ));
AOI21X2 U1754  (.A0 ( n1977 ) , .A1 ( n1965 ) , .B0 ( n1964 ) , .Y ( n1966 ));
NAND2BX4 U1755  (.AN ( n2082 ) , .B ( n2081 ) , .Y ( n2084 ));
INVX4 U1756  (.A ( n1852 ) , .Y ( n1871 ));
AOI21X2 U1757  (.A0 ( n2076 ) , .A1 ( n1948 ) , .B0 ( n1947 ) , .Y ( n1955 ));
INVX4 U1758  (.A ( n2014 ) , .Y ( n1965 ));
OAI21X1 U1759  (.A0 ( n2018 ) , .A1 ( n2002 ) , .B0 ( n1978 ) , .Y ( n1947 ));
AND2X4 U1760  (.A ( n1934 ) , .B ( n2018 ) , .Y ( n1936 ));
AOI21X6 U1761  (.A0 ( n1991 ) , .A1 ( n1996 ) , .B0 ( n1994 ) , .Y ( n1886 ));
NAND2X6 U1762  (.A ( n1664 ) , .B ( n1663 ) , .Y ( n1996 ));
NAND2X6 U1763  (.A ( n1776 ) , .B ( n1774 ) , .Y ( n2055 ));
NAND2X4 U1764  (.A ( n1859 ) , .B ( n1858 ) , .Y ( n1861 ));
NAND2BX4 U1765  (.AN ( n1776 ) , .B ( n1775 ) , .Y ( n2056 ));
XOR2X1 U1766  (.A ( n1946 ) , .B ( n2213 ) , .Y ( n1948 ));
NAND2X6 U1767  (.A ( n1604 ) , .B ( n1603 ) , .Y ( n1992 ));
NAND3X4 U1768  (.A ( n1676 ) , .B ( n1675 ) , .C ( n1674 ) , .Y ( n1704 ));
AOI21X1 U1769  (.A0 ( n2210 ) , .A1 ( n2108 ) , .B0 ( n2290 ) , .Y ( n1914 ));
NAND2X8 U1770  (.A ( n1755 ) , .B ( n1753 ) , .Y ( n1806 ));
NAND2X2 U1771  (.A ( n1930 ) , .B ( n1929 ) , .Y ( n1933 ));
XOR2X4 U1772  (.A ( n1590 ) , .B ( n1589 ) , .Y ( n1666 ));
OAI21X1 U1773  (.A0 ( n2017 ) , .A1 ( n2002 ) , .B0 ( n1978 ) , .Y ( n1913 ));
NAND2X4 U1774  (.A ( n1737 ) , .B ( n1729 ) , .Y ( n1740 ));
AND2X6 U1775  (.A ( n1608 ) , .B ( n1734 ) , .Y ( n1672 ));
AOI21X1 U1776  (.A0 ( n2107 ) , .A1 ( n2105 ) , .B0 ( n2290 ) , .Y ( n2109 ));
AND2X4 U1777  (.A ( n1644 ) , .B ( n1643 ) , .Y ( n1731 ));
NAND2X4 U1778  (.A ( n1499 ) , .B ( n1500 ) , .Y ( n1504 ));
NAND2X8 U1779  (.A ( n1588 ) , .B ( n1587 ) , .Y ( n1736 ));
NOR2BX1 U1780  (.AN ( n2097 ) , .B ( n2096 ) , .Y ( n2099 ));
AND2X6 U1781  (.A ( n1483 ) , .B ( n1482 ) , .Y ( n1499 ));
NAND2X6 U1782  (.A ( n1481 ) , .B ( n1480 ) , .Y ( n1500 ));
INVX1 U1783  (.A ( n2104 ) , .Y ( n2105 ));
INVX1 U1784  (.A ( n2095 ) , .Y ( n2096 ));
NAND2X4 U1785  (.A ( n1844 ) , .B ( n1843 ) , .Y ( n1864 ));
INVX4 U1786  (.A ( n1406 ) , .Y ( n1401 ));
AOI21XL U1787  (.A0 ( n2065 ) , .A1 ( n2064 ) , .B0 ( n2290 ) , .Y ( n2067 ));
OR2X6 U1788  (.A ( n1351 ) , .B ( n1350 ) , .Y ( n1506 ));
NAND3X6 U1789  (.A ( n1391 ) , .B ( n1390 ) , .C ( n1389 ) , .Y ( n1406 ));
INVX1 U1790  (.A ( n1387 ) , .Y ( n1221 ));
INVX4 U1791  (.A ( n1558 ) , .Y ( n1556 ));
INVXL U1792  (.A ( n2063 ) , .Y ( n2064 ));
CLKNAND2X2 U1793  (.A ( n1224 ) , .B ( n1223 ) , .Y ( n1226 ));
AND2X6 U1794  (.A ( n1816 ) , .B ( n1768 ) , .Y ( n1769 ));
NAND2X4 U1795  (.A ( n1055 ) , .B ( \intadd_7/SUM[1] ) , .Y ( n1558 ));
XOR2X1 U1796  (.A ( n1781 ) , .B ( n1779 ) , .Y ( n1754 ));
XOR2XL U1797  (.A ( n2052 ) , .B ( n2051 ) , .Y ( n2053 ));
OAI21X6 U1798  (.A0 ( n1455 ) , .A1 ( n1454 ) , .B0 ( n1453 ) , .Y ( n1516 ));
NAND2X2 U1799  (.A ( n1796 ) , .B ( n1795 ) , .Y ( n1813 ));
NAND2X6 U1800  (.A ( n1174 ) , .B ( n1173 ) , .Y ( n1340 ));
OAI21X4 U1801  (.A0 ( n1722 ) , .A1 ( n1721 ) , .B0 ( n1720 ) , .Y ( n1724 ));
XOR2XL U1802  (.A ( n1661 ) , .B ( n1720 ) , .Y ( n1662 ));
NAND2X4 U1803  (.A ( n1334 ) , .B ( n1333 ) , .Y ( n1335 ));
CLKXOR2X2 U1804  (.A ( n1719 ) , .B ( n1756 ) , .Y ( n1725 ));
NAND2X2 U1805  (.A ( n1625 ) , .B ( n1624 ) , .Y ( n1626 ));
OAI21X6 U1806  (.A0 ( n1157 ) , .A1 ( n1147 ) , .B0 ( n1146 ) , .Y ( n1168 ));
OAI21X1 U1807  (.A0 ( n1546 ) , .A1 ( n1545 ) , .B0 ( n1649 ) , .Y ( n1550 ));
XOR2X1 U1808  (.A ( n1464 ) , .B ( n1349 ) , .Y ( n1466 ));
OAI21X6 U1809  (.A0 ( n1294 ) , .A1 ( n1291 ) , .B0 ( n1292 ) , .Y ( n1286 ));
OAI21X6 U1810  (.A0 ( n1156 ) , .A1 ( n1145 ) , .B0 ( n1159 ) , .Y ( n1146 ));
XOR2X1 U1811  (.A ( n1679 ) , .B ( n1683 ) , .Y ( n1640 ));
OAI21X1 U1812  (.A0 ( n1464 ) , .A1 ( n1610 ) , .B0 ( n1463 ) , .Y ( n1465 ));
XOR2X1 U1813  (.A ( n1621 ) , .B ( n1622 ) , .Y ( n1584 ));
NAND2BX4 U1814  (.AN ( n1232 ) , .B ( n1210 ) , .Y ( n1214 ));
OAI2BB1X1 U1815  (.A0N ( n1716 ) , .A1N ( n1715 ) , .B0 ( n1763 ) , .Y ( n1717 ));
NAND2X4 U1816  (.A ( n2651 ) , .B ( n2556 ) , .Y ( n2296 ));
OAI21X2 U1817  (.A0 ( n1579 ) , .A1 ( n1578 ) , .B0 ( n1577 ) , .Y ( n1631 ));
XOR2X4 U1818  (.A ( n1163 ) , .B ( n1162 ) , .Y ( n1209 ));
OAI21X1 U1819  (.A0 ( n2698 ) , .A1 ( n1686 ) , .B0 ( n1611 ) , .Y ( n1612 ));
XOR2X1 U1820  (.A ( n1782 ) , .B ( n1784 ) , .Y ( n1752 ));
NAND2BX4 U1821  (.AN ( n1348 ) , .B ( n1347 ) , .Y ( n1463 ));
OAI21X6 U1822  (.A0 ( n1140 ) , .A1 ( n1139 ) , .B0 ( n1138 ) , .Y ( n1162 ));
NOR2BX1 U1823  (.AN ( n1306 ) , .B ( n1321 ) , .Y ( n1307 ));
BUFX10 U1824  (.A ( n1077 ) , .Y ( n1707 ));
NOR2X1 U1825  (.A ( n1202 ) , .B ( n1260 ) , .Y ( n1203 ));
MXI2X1 U1826  (.A ( n1848 ) , .B ( n1847 ) , .S0 ( n1866 ) , .Y ( n1849 ));
NOR2BX1 U1827  (.AN ( \intadd_4/n1  ) , .B ( n2289 ) , .Y ( n1912 ));
OAI21X1 U1828  (.A0 ( n1830 ) , .A1 ( n1049 ) , .B0 ( n2761 ) , .Y ( n1750 ));
XOR2X2 U1829  (.A ( n1161 ) , .B ( n1160 ) , .Y ( n1163 ));
OAI21X4 U1830  (.A0 ( n1234 ) , .A1 ( n1233 ) , .B0 ( n1235 ) , .Y ( n1138 ));
OAI21X1 U1831  (.A0 ( n1252 ) , .A1 ( n1472 ) , .B0 ( n1522 ) , .Y ( n1398 ));
NAND2X5 U1832  (.A ( n1137 ) , .B ( n1136 ) , .Y ( n1135 ));
AOI21X4 U1833  (.A0 ( n1170 ) , .A1 ( n1237 ) , .B0 ( n1128 ) , .Y ( n1116 ));
OAI21X1 U1834  (.A0 ( n1431 ) , .A1 ( n1430 ) , .B0 ( n1429 ) , .Y ( n1443 ));
XOR2X4 U1835  (.A ( n1123 ) , .B ( n1122 ) , .Y ( n1137 ));
BUFX10 U1836  (.A ( n1080 ) , .Y ( n2734 ));
MXI2X6 U1837  (.A ( n1072 ) , .B ( n1093 ) , .S0 ( n1071 ) , .Y ( n1073 ));
XOR2X2 U1838  (.A ( n1133 ) , .B ( n1132 ) , .Y ( n1238 ));
OAI21X2 U1839  (.A0 ( n2118 ) , .A1 ( n1802 ) , .B0 ( n1801 ) , .Y ( n1810 ));
XOR2X2 U1840  (.A ( n1110 ) , .B ( n1109 ) , .Y ( n1111 ));
NOR2BX1 U1841  (.AN ( n1492 ) , .B ( n2748 ) , .Y ( n1420 ));
AOI2BB1X1 U1842  (.A0N ( n1799 ) , .A1N ( n1430 ) , .B0 ( n1655 ) , .Y ( n1421 ));
BUFX10 U1843  (.A ( n1087 ) , .Y ( n1492 ));
INVX1 U1844  (.A ( n1628 ) , .Y ( n1630 ));
AND2X6 U1845  (.A ( n2556 ) , .B ( a[8] ) , .Y ( n1819 ));
NOR2BX1 U1846  (.AN ( b[6] ) , .B ( n1049 ) , .Y ( n1786 ));
NOR2BX1 U1847  (.AN ( n1119 ) , .B ( b[5] ) , .Y ( n1058 ));
NOR2X1 U1848  (.A ( \intadd_4/SUM[1] ) , .B ( n1949 ) , .Y ( n1918 ));
NOR2X1 U1849  (.A ( n1580 ) , .B ( n1049 ) , .Y ( n1581 ));
NOR2X1 U1850  (.A ( n2150 ) , .B ( c[12] ) , .Y ( n2155 ));
INVX1 U1851  (.A ( n1984 ) , .Y ( n1051 ));
INVX4 U1852  (.A ( n2749 ) , .Y ( n2655 ));
XOR2X1 U1853  (.A ( a[7] ) , .B ( b[7] ) , .Y ( n1246 ));
INVX4 U1854  (.A ( a[4] ) , .Y ( n1071 ));
NOR2X1 U1855  (.A ( c[11] ) , .B ( c[10] ) , .Y ( n2149 ));
NOR4X1 U1856  (.A ( b[7] ) , .B ( b[13] ) , .C ( b[11] ) , .D ( b[12] ) , .Y ( n1875 ));
NAND3BX4 U1857  (.AN ( clk ) , .B ( clk ) , .C ( clk ) , .Y ( n2608 ));
AOI222X4 U1858  (.A0 ( n2671 ) , .A1 ( n2636 ) , .B0 ( n2663 ) , .B1 ( n2659 ) , .C0 ( n2581 ) , .C1 ( n2305 ) , .Y ( n2712 ));
AOI21X4 U1859  (.A0 ( n1273 ) , .A1 ( n1231 ) , .B0 ( n1207 ) , .Y ( n1100 ));
NAND2X4 U1860  (.A ( n1100 ) , .B ( n1099 ) , .Y ( n1274 ));
MXI2X2 U1861  (.A ( n2232 ) , .B ( n2244 ) , .S0 ( n2241 ) , .Y ( n2279 ));
INVX4 U1862  (.A ( n1393 ) , .Y ( n1394 ));
NAND2X4 U1863  (.A ( n1325 ) , .B ( n1182 ) , .Y ( n1185 ));
NAND2X2 U1864  (.A ( n1502 ) , .B ( n1500 ) , .Y ( n1486 ));
AOI21X6 U1865  (.A0 ( n2094 ) , .A1 ( n2093 ) , .B0 ( n2092 ) , .Y ( n2134 ));
NAND2X2 U1866  (.A ( n1564 ) , .B ( n1563 ) , .Y ( n1565 ));
XOR2X8 U1867  (.A ( n1344 ) , .B ( n1331 ) , .Y ( n1377 ));
AOI21X4 U1868  (.A0 ( n2663 ) , .A1 ( n2671 ) , .B0 ( n2662 ) , .Y ( n2711 ));
OAI222X1 U1869  (.A0 ( n2658 ) , .A1 ( n2675 ) , .B0 ( n2674 ) , .B1 ( n2657 ) , .C0 ( n2678 ) , .C1 ( n2687 ) , .Y ( n2661 ));
AOI2BB2X4 U1870  (.B0 ( n2143 ) , .B1 ( n2181 ) , .A0N ( n2142 ) , .A1N ( n2141 ) , .Y ( n2144 ));
AND2X8 U1871  (.A ( n2514 ) , .B ( n2601 ) , .Y ( n2571 ));
NAND2BX4 U1872  (.AN ( n2211 ) , .B ( n2054 ) , .Y ( n2060 ));
NOR2BX4 U1873  (.AN ( n1569 ) , .B ( n1568 ) , .Y ( n1570 ));
AOI2BB2X4 U1874  (.B0 ( n2736 ) , .B1 ( n2517 ) , .A0N ( n2516 ) , .A1N ( n2515 ) , .Y ( n2535 ));
NOR2X4 U1875  (.A ( n1575 ) , .B ( n1176 ) , .Y ( n1353 ));
NAND3X4 U1876  (.A ( n2305 ) , .B ( n2374 ) , .C ( n2357 ) , .Y ( n2328 ));
XOR2X8 U1877  (.A ( n1336 ) , .B ( n1335 ) , .Y ( n1375 ));
XOR2X4 U1878  (.A ( n1486 ) , .B ( n1485 ) , .Y ( n1548 ));
INVX2 U1879  (.A ( n1300 ) , .Y ( n1304 ));
MXI2X6 U1880  (.A ( n2519 ) , .B ( n2548 ) , .S0 ( n2161 ) , .Y ( n2504 ));
MXI2X6 U1881  (.A ( n2522 ) , .B ( n2523 ) , .S0 ( n2189 ) , .Y ( n2601 ));
MXI2X4 U1882  (.A ( n2716 ) , .B ( n2646 ) , .S0 ( n2655 ) , .Y ( n1005 ));
NAND2X4 U1883  (.A ( n2198 ) , .B ( n2197 ) , .Y ( n2200 ));
NAND2BX4 U1884  (.AN ( n2469 ) , .B ( n2463 ) , .Y ( n2467 ));
NAND2BX8 U1885  (.AN ( n2353 ) , .B ( n2351 ) , .Y ( n2492 ));
AOI211X4 U1886  (.A0 ( n2547 ) , .A1 ( n2305 ) , .B0 ( n2546 ) , .C0 ( n2545 ) , .Y ( n2713 ));
XOR2X4 U1887  (.A ( n1411 ) , .B ( n1410 ) , .Y ( n1415 ));
XOR2X8 U1888  (.A ( n1926 ) , .B ( n1925 ) , .Y ( n2007 ));
NAND2X8 U1889  (.A ( n1859 ) , .B ( n1837 ) , .Y ( n2081 ));
XNOR2X4 U1890  (.A ( n1516 ) , .B ( n1462 ) , .Y ( n1468 ));
OR2X6 U1891  (.A ( n2475 ) , .B ( n2476 ) , .Y ( n2478 ));
XOR2X8 U1892  (.A ( n1646 ) , .B ( n1645 ) , .Y ( n1668 ));
NAND2X4 U1893  (.A ( n1736 ) , .B ( n1607 ) , .Y ( n1608 ));
OAI211X4 U1894  (.A0 ( n2505 ) , .A1 ( c[10] ) , .B0 ( n2138 ) , .C0 ( n2140 ) , .Y ( n1986 ));
AOI22X2 U1895  (.A0 ( n2639 ) , .A1 ( n2690 ) , .B0 ( n2689 ) , .B1 ( n2638 ) , .Y ( n2640 ));
OAI21X2 U1896  (.A0 ( n2642 ) , .A1 ( n2641 ) , .B0 ( n2640 ) , .Y ( n2645 ));
NAND2BX8 U1897  (.AN ( n1357 ) , .B ( n1361 ) , .Y ( n1369 ));
CLKBUFX40 U1898  (.A ( n2161 ) , .Y ( n2189 ));
NAND3X4 U1899  (.A ( n1495 ) , .B ( n1494 ) , .C ( n1493 ) , .Y ( n1599 ));
NAND2X2 U1900  (.A ( n1563 ) , .B ( n1555 ) , .Y ( n1560 ));
AOI211X2 U1901  (.A0 ( n2684 ) , .A1 ( n2670 ) , .B0 ( n2649 ) , .C0 ( n2648 ) , .Y ( n2652 ));
OAI22X1 U1902  (.A0 ( n2687 ) , .A1 ( n2675 ) , .B0 ( n2674 ) , .B1 ( n2679 ) , .Y ( n2649 ));
AOI22X4 U1903  (.A0 ( n2671 ) , .A1 ( n2654 ) , .B0 ( n2556 ) , .B1 ( n2653 ) , .Y ( n2717 ));
AOI21X8 U1904  (.A0 ( n2168 ) , .A1 ( n2166 ) , .B0 ( n2165 ) , .Y ( n2175 ));
OAI22X4 U1905  (.A0 ( n2607 ) , .A1 ( n2606 ) , .B0 ( n2605 ) , .B1 ( n2722 ) , .Y ( n999 ));
OAI21X8 U1906  (.A0 ( n1371 ) , .A1 ( n1370 ) , .B0 ( n1346 ) , .Y ( n1467 ));
OA21X4 U1907  (.A0 ( n1371 ) , .A1 ( n1369 ) , .B0 ( n1345 ) , .Y ( n1346 ));
NAND2X2 U1908  (.A ( n1484 ) , .B ( n1501 ) , .Y ( n1485 ));
NAND2BX4 U1909  (.AN ( n2111 ) , .B ( n2110 ) , .Y ( n2113 ));
NAND2BX8 U1910  (.AN ( n1352 ) , .B ( n1351 ) , .Y ( n1507 ));
AND4X4 U1911  (.A ( n2536 ) , .B ( n2535 ) , .C ( n2534 ) , .D ( n1050 ) , .Y ( n2609 ));
OAI21X4 U1912  (.A0 ( n1567 ) , .A1 ( n1566 ) , .B0 ( n1565 ) , .Y ( n1572 ));
NOR2X6 U1913  (.A ( n2642 ) , .B ( n2600 ) , .Y ( n2570 ));
NAND3X2 U1914  (.A ( n1121 ) , .B ( n1427 ) , .C ( n2020 ) , .Y ( n1132 ));
NAND2X2 U1915  (.A ( n1285 ) , .B ( n1284 ) , .Y ( n1287 ));
BUFX8 U1916  (.A ( n1111 ) , .Y ( n1582 ));
AND2X4 U1917  (.A ( n1728 ) , .B ( n1674 ) , .Y ( n1645 ));
AOI21X4 U1918  (.A0 ( n1670 ) , .A1 ( n1605 ) , .B0 ( n1607 ) , .Y ( n1590 ));
OAI21XL U1919  (.A0 ( n1655 ) , .A1 ( n1430 ) , .B0 ( n1428 ) , .Y ( n1429 ));
NAND2BXL U1920  (.AN ( n2556 ) , .B ( c[2] ) , .Y ( n2335 ));
NAND2BXL U1921  (.AN ( n2556 ) , .B ( c[4] ) , .Y ( n2310 ));
AND2X2 U1922  (.A ( n1374 ) , .B ( n1358 ) , .Y ( n1356 ));
OR2X4 U1923  (.A ( n1338 ) , .B ( n1340 ) , .Y ( n1337 ));
NAND2X2 U1924  (.A ( n1492 ) , .B ( n1121 ) , .Y ( n1122 ));
AOI21X4 U1925  (.A0 ( n1133 ) , .A1 ( n2020 ) , .B0 ( n1239 ) , .Y ( n1136 ));
NAND2X2 U1926  (.A ( n1506 ) , .B ( n1561 ) , .Y ( n1451 ));
OAI21X4 U1927  (.A0 ( n1842 ) , .A1 ( n1841 ) , .B0 ( n1840 ) , .Y ( n1844 ));
NAND2X4 U1928  (.A ( n1887 ) , .B ( n2042 ) , .Y ( n1893 ));
NAND3X4 U1929  (.A ( n2042 ) , .B ( n1993 ) , .C ( n1890 ) , .Y ( n1892 ));
MXI2XL U1930  (.A ( n1976 ) , .B ( n1975 ) , .S0 ( n1974 ) , .Y ( n1981 ));
OAI211X2 U1931  (.A0 ( n2679 ) , .A1 ( n2633 ) , .B0 ( n2498 ) , .C0 ( n2497 ) , .Y ( n2499 ));
NAND2X8 U1932  (.A ( n2583 ) , .B ( n2459 ) , .Y ( n2686 ));
AND2X2 U1933  (.A ( n2676 ) , .B ( n2673 ) , .Y ( n2459 ));
OAI21X2 U1934  (.A0 ( n1304 ) , .A1 ( n1303 ) , .B0 ( n1302 ) , .Y ( n1332 ));
NAND2X2 U1935  (.A ( n1308 ) , .B ( n1309 ) , .Y ( n1333 ));
NAND2X2 U1936  (.A ( n1297 ) , .B ( n1296 ) , .Y ( n1366 ));
AND2X2 U1937  (.A ( n1169 ) , .B ( n1117 ) , .Y ( n1145 ));
CLKXOR2X2 U1938  (.A ( n1467 ) , .B ( n1466 ) , .Y ( n1350 ));
OA21X2 U1939  (.A0 ( n1100 ) , .A1 ( n1099 ) , .B0 ( n1274 ) , .Y ( n1103 ));
AOI21X4 U1940  (.A0 ( n1364 ) , .A1 ( n1363 ) , .B0 ( n1362 ) , .Y ( n1393 ));
OAI21X1 U1941  (.A0 ( n1361 ) , .A1 ( n1375 ) , .B0 ( n1379 ) , .Y ( n1362 ));
NAND2X4 U1942  (.A ( n1510 ) , .B ( n1506 ) , .Y ( n1567 ));
NAND2X4 U1943  (.A ( b[7] ) , .B ( n2556 ) , .Y ( n1686 ));
INVX4 U1944  (.A ( n1145 ) , .Y ( n1157 ));
INVX2 U1945  (.A ( n1450 ) , .Y ( n1561 ));
CLKXOR2X4 U1946  (.A ( n1693 ) , .B ( n1619 ) , .Y ( n1641 ));
XOR2X1 U1947  (.A ( n1594 ) , .B ( n1593 ) , .Y ( n1544 ));
XOR2XL U1948  (.A ( n1865 ) , .B ( n1049 ) , .Y ( n1847 ));
INVX2 U1949  (.A ( n1208 ) , .Y ( n1182 ));
NAND2X2 U1950  (.A ( n1490 ) , .B ( n1489 ) , .Y ( n1491 ));
NOR2X6 U1951  (.A ( n1669 ) , .B ( n1606 ) , .Y ( n1729 ));
CLKXOR2X2 U1952  (.A ( n1127 ) , .B ( n1135 ) , .Y ( n1161 ));
NAND2X2 U1953  (.A ( n1134 ) , .B ( n1238 ) , .Y ( n1234 ));
OR2X4 U1954  (.A ( a[1] ) , .B ( \u_mac/mul/N7  ) , .Y ( n1084 ));
AND2X2 U1955  (.A ( n1427 ) , .B ( n1657 ) , .Y ( n1489 ));
INVX2 U1956  (.A ( n1733 ) , .Y ( n1607 ));
INVX2 U1957  (.A ( n1588 ) , .Y ( n1586 ));
INVXL U1958  (.A ( n2117 ) , .Y ( n2120 ));
NAND2X4 U1959  (.A ( n1209 ) , .B ( n1208 ) , .Y ( n1212 ));
NAND2X4 U1960  (.A ( n1549 ) , .B ( n1550 ) , .Y ( n1924 ));
NAND2XL U1961  (.A ( n1121 ) , .B ( n1819 ) , .Y ( n1414 ));
INVX4 U1962  (.A ( \u_mac/mul/N7  ) , .Y ( n1430 ));
OAI22XL U1963  (.A0 ( n2016 ) , .A1 ( c[1] ) , .B0 ( n2018 ) , .B1 ( c[0] ) , .Y ( n2024 ));
INVXL U1964  (.A ( n1536 ) , .Y ( n1497 ));
XOR2XL U1965  (.A ( n1988 ) , .B ( n1987 ) , .Y ( n1990 ));
NAND2BX2 U1966  (.AN ( n2177 ) , .B ( n2176 ) , .Y ( n2178 ));
NAND2XL U1967  (.A ( n1241 ) , .B ( n1240 ) , .Y ( n2004 ));
XOR2XL U1968  (.A ( n1910 ) , .B ( n2066 ) , .Y ( n1248 ));
NAND2BX4 U1969  (.AN ( n2152 ) , .B ( c[12] ) , .Y ( n2135 ));
NAND3X4 U1970  (.A ( n2040 ) , .B ( n2042 ) , .C ( n2055 ) , .Y ( n1778 ));
OAI21X4 U1971  (.A0 ( n2083 ) , .A1 ( n2111 ) , .B0 ( n1869 ) , .Y ( n1870 ));
INVX2 U1972  (.A ( n2234 ) , .Y ( n2201 ));
AND2X2 U1973  (.A ( n1548 ) , .B ( n1547 ) , .Y ( n1928 ));
AOI21XL U1974  (.A0 ( n2037 ) , .A1 ( n2036 ) , .B0 ( n2290 ) , .Y ( n2038 ));
NAND3X4 U1975  (.A ( n2073 ) , .B ( n2072 ) , .C ( n2071 ) , .Y ( n2382 ));
NAND2X4 U1976  (.A ( n2340 ) , .B ( n2339 ) , .Y ( n2332 ));
NAND2BXL U1977  (.AN ( n2556 ) , .B ( c[7] ) , .Y ( n2390 ));
INVXL U1978  (.A ( n2390 ) , .Y ( n2391 ));
AND2X2 U1979  (.A ( n2455 ) , .B ( n2485 ) , .Y ( n2401 ));
OAI21X1 U1980  (.A0 ( n1965 ) , .A1 ( n2002 ) , .B0 ( n1978 ) , .Y ( n1964 ));
NOR2XL U1981  (.A ( n1976 ) , .B ( n1973 ) , .Y ( n1975 ));
OAI21XL U1982  (.A0 ( n1951 ) , .A1 ( \intadd_4/SUM[0] ) , .B0 ( n1950 ) , .Y ( n1952 ));
AND2X2 U1983  (.A ( n1246 ) , .B ( n2692 ) , .Y ( n2076 ));
NAND2X4 U1984  (.A ( n2464 ) , .B ( n2465 ) , .Y ( n2438 ));
NAND2BXL U1985  (.AN ( n2214 ) , .B ( n2213 ) , .Y ( n2215 ));
NAND2BXL U1986  (.AN ( n2211 ) , .B ( n2210 ) , .Y ( n2217 ));
AND2X2 U1987  (.A ( n2332 ) , .B ( n2305 ) , .Y ( n2338 ));
INVXL U1988  (.A ( n2674 ) , .Y ( n2489 ));
INVX2 U1989  (.A ( n2076 ) , .Y ( n2290 ));
NOR2XL U1990  (.A ( n2523 ) , .B ( n2556 ) , .Y ( n2524 ));
INVX2 U1991  (.A ( n2152 ) , .Y ( n2522 ));
MXI2X4 U1992  (.A ( n2345 ) , .B ( c[0] ) , .S0 ( n2692 ) , .Y ( n2475 ));
XOR2XL U1993  (.A ( b[15] ) , .B ( a[15] ) , .Y ( n2288 ));
XOR2X1 U1994  (.A ( n2623 ) , .B ( n2595 ) , .Y ( n2538 ));
XNOR2XL U1995  (.A ( n2595 ) , .B ( n2627 ) , .Y ( n2544 ));
XOR2XL U1996  (.A ( n2540 ) , .B ( c[11] ) , .Y ( n2541 ));
OAI22XL U1997  (.A0 ( n2680 ) , .A1 ( n2679 ) , .B0 ( n2678 ) , .B1 ( n2677 ) , .Y ( n2681 ));
INVX2 U1998  (.A ( n2651 ) , .Y ( n2690 ));
INVXL U1999  (.A ( n2517 ) , .Y ( n2515 ));
INVXL U2000  (.A ( n2592 ) , .Y ( n2526 ));
NAND2XL U2001  (.A ( n2531 ) , .B ( n2552 ) , .Y ( n2532 ));
INVXL U2002  (.A ( n2553 ) , .Y ( n2531 ));
CLKXOR2X2 U2003  (.A ( n2292 ) , .B ( n2291 ) , .Y ( n2651 ));
AOI21X4 U2004  (.A0 ( n2456 ) , .A1 ( n2458 ) , .B0 ( n2427 ) , .Y ( n2431 ));
AND2X2 U2005  (.A ( \intadd_4/SUM[2] ) , .B ( n1957 ) , .Y ( n1960 ));
INVXL U2006  (.A ( c[7] ) , .Y ( n2503 ));
AND2X2 U2007  (.A ( n2671 ) , .B ( n2638 ) , .Y ( n1053 ));
INVXL U2008  (.A ( n2627 ) , .Y ( n2626 ));
NAND2XL U2009  (.A ( n2593 ) , .B ( n2592 ) , .Y ( n2594 ));
AOI21XL U2010  (.A0 ( n2595 ) , .A1 ( n2627 ) , .B0 ( n2601 ) , .Y ( n2596 ));
NOR3X2 U2011  (.A ( n2571 ) , .B ( n2570 ) , .C ( n2569 ) , .Y ( n2573 ));
XOR2X1 U2012  (.A ( n2560 ) , .B ( n2559 ) , .Y ( n2745 ));
NAND2XL U2013  (.A ( n2613 ) , .B ( n2611 ) , .Y ( n2559 ));
INVXL U2014  (.A ( c[2] ) , .Y ( n2582 ));
MXI2X4 U2015  (.A ( n2609 ) , .B ( n2537 ) , .S0 ( n2655 ) , .Y ( n998 ));
NOR2XL U2016  (.A ( c[12] ) , .B ( n2749 ) , .Y ( n2606 ));
INVXL U2017  (.A ( n2599 ) , .Y ( n2605 ));
MX2XL U2018  (.A ( b[1] ) , .B ( in_b[1] ) , .S0 ( n2749 ) , .Y ( n1030 ));
MXI2X1 U2019  (.A ( n2712 ) , .B ( n2582 ) , .S0 ( n2655 ) , .Y ( n1009 ));
MX2XL U2020  (.A ( b[7] ) , .B ( in_b[7] ) , .S0 ( n2749 ) , .Y ( n1036 ));
NAND2X2 U2021  (.A ( n1540 ) , .B ( n1539 ) , .Y ( n1537 ));
NAND2BX4 U2022  (.AN ( n2211 ) , .B ( n2039 ) , .Y ( n2046 ));
NOR2X8 U2023  (.A ( n1895 ) , .B ( n1852 ) , .Y ( n2115 ));
XOR2X8 U2024  (.A ( n1471 ) , .B ( n1470 ) , .Y ( n1481 ));
NAND3X4 U2025  (.A ( n1452 ) , .B ( n1451 ) , .C ( n1507 ) , .Y ( n1471 ));
NAND4X4 U2026  (.A ( n2509 ) , .B ( n2678 ) , .C ( n2680 ) , .D ( n2674 ) , .Y ( n2513 ));
AOI21X4 U2027  (.A0 ( n2413 ) , .A1 ( n2412 ) , .B0 ( n2550 ) , .Y ( n2414 ));
XNOR2X2 U2028  (.A ( n1368 ) , .B ( n1367 ) , .Y ( n1385 ));
CLKXOR2X8 U2029  (.A ( n1120 ) , .B ( b[1] ) , .Y ( n1121 ));
XOR2X1 U2030  (.A ( a[10] ) , .B ( b[10] ) , .Y ( n1951 ));
MXI2X1 U2031  (.A ( n2720 ) , .B ( n2483 ) , .S0 ( n2655 ) , .Y ( n1011 ));
INVX2 U2032  (.A ( c[6] ) , .Y ( n2646 ));
NAND2BXL U2033  (.AN ( n2556 ) , .B ( c[6] ) , .Y ( n2380 ));
NOR4XL U2034  (.A ( b[8] ) , .B ( b[9] ) , .C ( b[14] ) , .D ( b[15] ) , .Y ( n1874 ));
NOR4XL U2035  (.A ( a[8] ) , .B ( a[9] ) , .C ( a[14] ) , .D ( a[15] ) , .Y ( n1879 ));
NOR4XL U2036  (.A ( a[6] ) , .B ( a[13] ) , .C ( a[11] ) , .D ( a[12] ) , .Y ( n1880 ));
INVXL U2037  (.A ( c[1] ) , .Y ( n2672 ));
NAND3XL U2038  (.A ( n2224 ) , .B ( n2223 ) , .C ( n2222 ) , .Y ( n2348 ));
OAI2BB1X2 U2039  (.A0N ( n1406 ) , .A1N ( n1405 ) , .B0 ( n1404 ) , .Y ( n1411 ));
NAND3X4 U2040  (.A ( n1409 ) , .B ( n1406 ) , .C ( n1405 ) , .Y ( n1450 ));
AO21X4 U2041  (.A0 ( n1516 ) , .A1 ( n1515 ) , .B0 ( n1514 ) , .Y ( n1055 ));
AO21X4 U2042  (.A0 ( n1286 ) , .A1 ( n1285 ) , .B0 ( n1277 ) , .Y ( n1056 ));
INVXL U2043  (.A ( c[8] ) , .Y ( n2131 ));
INVX2 U2044  (.A ( n1284 ) , .Y ( n1277 ));
CLKXOR2X2 U2045  (.A ( n1098 ) , .B ( n1097 ) , .Y ( n1099 ));
INVXL U2046  (.A ( n2020 ) , .Y ( n2003 ));
NAND2XL U2047  (.A ( n2013 ) , .B ( n2010 ) , .Y ( n2011 ));
INVXL U2048  (.A ( n1972 ) , .Y ( n1973 ));
NOR2XL U2049  (.A ( n2537 ) , .B ( n2556 ) , .Y ( n2529 ));
OR2X4 U2050  (.A ( b[1] ) , .B ( \u_mac/mul/N17  ) , .Y ( n1112 ));
NAND2BX8 U2051  (.AN ( n2293 ) , .B ( b[7] ) , .Y ( n1119 ));
NOR2X2 U2052  (.A ( n1119 ) , .B ( n1061 ) , .Y ( n1059 ));
INVX4 U2053  (.A ( a[2] ) , .Y ( n1085 ));
NAND2X8 U2054  (.A ( n1065 ) , .B ( n2760 ) , .Y ( n1095 ));
NAND2X8 U2055  (.A ( n1066 ) , .B ( n1071 ) , .Y ( n1074 ));
NAND2X2 U2056  (.A ( n1074 ) , .B ( n1093 ) , .Y ( n1067 ));
INVX4 U2057  (.A ( a[5] ) , .Y ( n1759 ));
NAND2BX2 U2058  (.AN ( n1091 ) , .B ( n2733 ) , .Y ( n2697 ));
NAND2BX8 U2059  (.AN ( n1073 ) , .B ( n1074 ) , .Y ( n1176 ));
NAND2X2 U2060  (.A ( n1707 ) , .B ( n2699 ) , .Y ( n2706 ));
NAND2X2 U2061  (.A ( n1877 ) , .B ( n1107 ) , .Y ( n1079 ));
XOR2X2 U2062  (.A ( n1079 ) , .B ( n2761 ) , .Y ( n1080 ));
NAND2X2 U2063  (.A ( n2734 ) , .B ( n2732 ) , .Y ( n2754 ));
AND2X2 U2064  (.A ( \intadd_4/SUM[0] ) , .B ( n1951 ) , .Y ( n1949 ));
AND2X2 U2065  (.A ( \intadd_4/SUM[1] ) , .B ( n1949 ) , .Y ( n1957 ));
CLKXOR2X2 U2066  (.A ( \intadd_4/SUM[3] ) , .B ( n1960 ) , .Y ( n1974 ));
NAND2BX4 U2067  (.AN ( n1088 ) , .B ( n1084 ) , .Y ( n1086 ));
NAND2X2 U2068  (.A ( n2699 ) , .B ( n1492 ) , .Y ( n1273 ));
NAND2X2 U2069  (.A ( n2699 ) , .B ( n2748 ) , .Y ( n1231 ));
BUFX5 U2070  (.A ( n1090 ) , .Y ( n1427 ));
NAND2BX2 U2071  (.AN ( n1091 ) , .B ( n1427 ) , .Y ( n1207 ));
INVX2 U2072  (.A ( n1492 ) , .Y ( n1487 ));
NAND2X2 U2073  (.A ( n1093 ) , .B ( n1092 ) , .Y ( n1094 ));
NAND2BX8 U2074  (.AN ( n1096 ) , .B ( n1095 ) , .Y ( n1118 ));
NOR2X2 U2075  (.A ( n1575 ) , .B ( n1118 ) , .Y ( n1097 ));
NAND2X2 U2076  (.A ( n2734 ) , .B ( n1427 ) , .Y ( n1269 ));
INVX4 U2077  (.A ( n1686 ) , .Y ( n2731 ));
OR2X2 U2078  (.A ( n1103 ) , .B ( n1102 ) , .Y ( n1256 ));
NAND2X2 U2079  (.A ( n1103 ) , .B ( n1102 ) , .Y ( n1253 ));
NAND2BX2 U2080  (.AN ( n1207 ) , .B ( n1231 ) , .Y ( n1104 ));
XOR2X1 U2081  (.A ( n1104 ) , .B ( n1273 ) , .Y ( n1202 ));
AND2X2 U2082  (.A ( n2734 ) , .B ( n2748 ) , .Y ( n1260 ));
AND2X2 U2083  (.A ( n1202 ) , .B ( n1260 ) , .Y ( n1255 ));
XNOR2X1 U2084  (.A ( n1105 ) , .B ( n1255 ) , .Y ( n1196 ));
INVX2 U2085  (.A ( n1106 ) , .Y ( n1108 ));
NAND2BX2 U2086  (.AN ( n1118 ) , .B ( n1582 ) , .Y ( n1172 ));
XOR2X8 U2087  (.A ( n1113 ) , .B ( n1580 ) , .Y ( n1315 ));
AND2X2 U2088  (.A ( n1315 ) , .B ( n1492 ) , .Y ( n1148 ));
INVX2 U2089  (.A ( n1315 ) , .Y ( n1474 ));
INVX2 U2090  (.A ( n1582 ) , .Y ( n1175 ));
OAI22X1 U2091  (.A0 ( n1118 ) , .A1 ( n1474 ) , .B0 ( n1487 ) , .B1 ( n1175 ) , .Y ( n1114 ));
AND2X2 U2092  (.A ( n1315 ) , .B ( n2748 ) , .Y ( n1134 ));
INVX2 U2093  (.A ( n1134 ) , .Y ( n1237 ));
NAND2X2 U2094  (.A ( n1582 ) , .B ( n1427 ) , .Y ( n1128 ));
NAND2BX8 U2095  (.AN ( n1115 ) , .B ( n1116 ) , .Y ( n1169 ));
NAND2BX2 U2096  (.AN ( n1116 ) , .B ( n1115 ) , .Y ( n1117 ));
NAND2BX2 U2097  (.AN ( n1118 ) , .B ( n2750 ) , .Y ( n1123 ));
INVX4 U2098  (.A ( n2750 ) , .Y ( n1403 ));
NAND2X4 U2099  (.A ( n1492 ) , .B ( n2750 ) , .Y ( n1133 ));
NAND2X2 U2100  (.A ( n2750 ) , .B ( n2748 ) , .Y ( n2020 ));
NAND2X2 U2101  (.A ( n1121 ) , .B ( n1427 ) , .Y ( n1239 ));
INVX2 U2102  (.A ( n1121 ) , .Y ( n1164 ));
NOR2X2 U2103  (.A ( n1118 ) , .B ( n1164 ) , .Y ( n1126 ));
INVX2 U2104  (.A ( n1126 ) , .Y ( n1124 ));
NAND2BX2 U2105  (.AN ( n1128 ) , .B ( n1237 ) , .Y ( n1125 ));
NAND2X2 U2106  (.A ( n1126 ) , .B ( n1133 ) , .Y ( n1127 ));
NAND2BX2 U2107  (.AN ( n1128 ) , .B ( n1134 ) , .Y ( n1131 ));
INVX2 U2108  (.A ( n1427 ) , .Y ( n1259 ));
NAND2X2 U2109  (.A ( n1582 ) , .B ( n2748 ) , .Y ( n1129 ));
OAI21X1 U2110  (.A0 ( n1259 ) , .A1 ( n1474 ) , .B0 ( n1129 ) , .Y ( n1130 ));
NAND2X2 U2111  (.A ( n1131 ) , .B ( n1130 ) , .Y ( n1233 ));
INVX2 U2112  (.A ( n1233 ) , .Y ( n1140 ));
INVX2 U2113  (.A ( n1234 ) , .Y ( n1139 ));
OAI21X1 U2114  (.A0 ( n1137 ) , .A1 ( n1136 ) , .B0 ( n1135 ) , .Y ( n1235 ));
NAND2X2 U2115  (.A ( n1161 ) , .B ( n1142 ) , .Y ( n1143 ));
XOR2X1 U2116  (.A ( n1169 ) , .B ( n1149 ) , .Y ( n1150 ));
XOR2X8 U2117  (.A ( n1168 ) , .B ( n1150 ) , .Y ( n1166 ));
NAND2BX2 U2118  (.AN ( n1176 ) , .B ( n1315 ) , .Y ( n1306 ));
NOR2X2 U2119  (.A ( n1176 ) , .B ( n1403 ) , .Y ( n1208 ));
NAND2X2 U2120  (.A ( n2733 ) , .B ( n1121 ) , .Y ( n1183 ));
NOR2BX4 U2121  (.AN ( n1182 ) , .B ( n1183 ) , .Y ( n1151 ));
NAND2X4 U2122  (.A ( n1707 ) , .B ( n2750 ) , .Y ( n1325 ));
XOR2X8 U2123  (.A ( n1151 ) , .B ( n1325 ) , .Y ( n1152 ));
INVX2 U2124  (.A ( n1306 ) , .Y ( n1153 ));
NAND2X2 U2125  (.A ( n1155 ) , .B ( n1181 ) , .Y ( n1198 ));
NAND2X2 U2126  (.A ( n1166 ) , .B ( n1198 ) , .Y ( n1359 ));
OAI22X1 U2127  (.A0 ( n1706 ) , .A1 ( n1164 ) , .B0 ( n1403 ) , .B1 ( n1177 ) , .Y ( n1165 ));
OAI21X1 U2128  (.A0 ( n1183 ) , .A1 ( n1182 ) , .B0 ( n1165 ) , .Y ( n1211 ));
NAND3X4 U2129  (.A ( n1171 ) , .B ( n1170 ) , .C ( n1169 ) , .Y ( n1174 ));
INVX2 U2130  (.A ( n1172 ) , .Y ( n1173 ));
NAND2X2 U2131  (.A ( n2733 ) , .B ( n1582 ) , .Y ( n1321 ));
OR2X2 U2132  (.A ( n1321 ) , .B ( n1306 ) , .Y ( n1319 ));
INVX2 U2133  (.A ( n1183 ) , .Y ( n1184 ));
NAND2X2 U2134  (.A ( n1185 ) , .B ( n1184 ) , .Y ( n1189 ));
AND2X6 U2135  (.A ( a[7] ) , .B ( n2556 ) , .Y ( n2702 ));
INVX2 U2136  (.A ( n1188 ) , .Y ( n1190 ));
NAND2X2 U2137  (.A ( n1190 ) , .B ( n1189 ) , .Y ( n1191 ));
OR2X4 U2138  (.A ( n1196 ) , .B ( n1195 ) , .Y ( n1388 ));
INVX2 U2139  (.A ( n1195 ) , .Y ( n1197 ));
NAND2BX4 U2140  (.AN ( n1197 ) , .B ( n1196 ) , .Y ( n1389 ));
INVX2 U2141  (.A ( n1220 ) , .Y ( n1205 ));
NAND2X2 U2142  (.A ( n1205 ) , .B ( n1204 ) , .Y ( n1223 ));
OAI22X1 U2143  (.A0 ( n1091 ) , .A1 ( n1430 ) , .B0 ( n1575 ) , .B1 ( n1259 ) , .Y ( n1206 ));
OAI21X1 U2144  (.A0 ( n1207 ) , .A1 ( n1231 ) , .B0 ( n1206 ) , .Y ( n1229 ));
ADDFHX4 U2145  (.A ( n1213 ) , .B ( n1212 ) , .CI ( n1211 ) , .CO ( n1201 ) , .S ( n1215 ));
NAND2X2 U2146  (.A ( n1214 ) , .B ( n1215 ) , .Y ( n1228 ));
NAND2BX2 U2147  (.AN ( n1229 ) , .B ( n1228 ) , .Y ( n1218 ));
INVX2 U2148  (.A ( n1215 ) , .Y ( n1216 ));
NAND2X2 U2149  (.A ( n1217 ) , .B ( n1216 ) , .Y ( n1227 ));
AND2X2 U2150  (.A ( n1220 ) , .B ( n1219 ) , .Y ( n1386 ));
INVX2 U2151  (.A ( n1386 ) , .Y ( n1224 ));
XOR2X1 U2152  (.A ( n1222 ) , .B ( n1052 ) , .Y ( n1910 ));
XOR2X1 U2153  (.A ( n1226 ) , .B ( n1225 ) , .Y ( n2062 ));
XOR2X1 U2154  (.A ( n1230 ) , .B ( n1229 ) , .Y ( n2052 ));
INVX2 U2155  (.A ( n2052 ) , .Y ( n1245 ));
XOR2X1 U2156  (.A ( n1232 ) , .B ( n1231 ) , .Y ( n2037 ));
XOR2X1 U2157  (.A ( n1236 ) , .B ( n1235 ) , .Y ( n1988 ));
XOR2X1 U2158  (.A ( n1238 ) , .B ( n1237 ) , .Y ( n2008 ));
NAND2BXL U2159  (.AN ( n1239 ) , .B ( n2003 ) , .Y ( n1241 ));
AO22XL U2160  (.A0 ( n2750 ) , .A1 ( n1427 ) , .B0 ( n2748 ) , .B1 ( n1121 ) , .Y ( n1240 ));
NAND2X2 U2161  (.A ( n1988 ) , .B ( n1987 ) , .Y ( n2036 ));
NAND2X2 U2162  (.A ( n1243 ) , .B ( n1242 ) , .Y ( n2051 ));
AND2X2 U2163  (.A ( n1245 ) , .B ( n1244 ) , .Y ( n2063 ));
NAND2X2 U2164  (.A ( n2062 ) , .B ( n2063 ) , .Y ( n2066 ));
AND2X2 U2165  (.A ( n1247 ) , .B ( n2692 ) , .Y ( n2106 ));
AOI22XL U2166  (.A0 ( n1248 ) , .A1 ( n2076 ) , .B0 ( n2106 ) , .B1 ( n1910 ) , .Y ( n1905 ));
AOI21X1 U2167  (.A0 ( n1412 ) , .A1 ( n1819 ) , .B0 ( n1049 ) , .Y ( n1249 ));
NAND2X2 U2168  (.A ( n1249 ) , .B ( n1121 ) , .Y ( n1250 ));
AND2X2 U2169  (.A ( n1315 ) , .B ( n1819 ) , .Y ( n1472 ));
INVX2 U2170  (.A ( n1253 ) , .Y ( n1254 ));
NAND2BX2 U2171  (.AN ( n1091 ) , .B ( n1264 ) , .Y ( n1272 ));
XNOR2X2 U2172  (.A ( n1274 ) , .B ( n1258 ) , .Y ( n1263 ));
NAND2X2 U2173  (.A ( n2734 ) , .B ( n1492 ) , .Y ( n1267 ));
XOR2X1 U2174  (.A ( n1261 ) , .B ( n1458 ) , .Y ( n1262 ));
NAND2X4 U2175  (.A ( n1263 ) , .B ( n1262 ) , .Y ( n1292 ));
NAND2X2 U2176  (.A ( n2734 ) , .B ( n1264 ) , .Y ( n1265 ));
OAI21X1 U2177  (.A0 ( n1686 ) , .A1 ( n1487 ) , .B0 ( n1265 ) , .Y ( n1266 ));
OA21X4 U2178  (.A0 ( n1456 ) , .A1 ( n1267 ) , .B0 ( n1266 ) , .Y ( n1271 ));
NOR2X2 U2179  (.A ( n1269 ) , .B ( n1268 ) , .Y ( n1270 ));
AND2X2 U2180  (.A ( n1271 ) , .B ( n1270 ) , .Y ( n1459 ));
AOI2BB1X2 U2181  (.A0N ( n1271 ) , .A1N ( n1270 ) , .B0 ( n1459 ) , .Y ( n1276 ));
OR2X2 U2182  (.A ( n1276 ) , .B ( n1275 ) , .Y ( n1285 ));
NAND2X2 U2183  (.A ( n1276 ) , .B ( n1275 ) , .Y ( n1284 ));
XOR2X1 U2184  (.A ( n1459 ) , .B ( n1278 ) , .Y ( n1279 ));
NOR2X4 U2185  (.A ( n1282 ) , .B ( n1281 ) , .Y ( n1455 ));
NAND2X2 U2186  (.A ( n1282 ) , .B ( n1281 ) , .Y ( n1453 ));
XNOR2X4 U2187  (.A ( n1287 ) , .B ( n1286 ) , .Y ( n1297 ));
AOI22XL U2188  (.A0 ( n1289 ) , .A1 ( n2732 ) , .B0 ( n2733 ) , .B1 ( n2699 ) , .Y ( n1290 ));
NOR2X2 U2189  (.A ( n2696 ) , .B ( n1290 ) , .Y ( n1296 ));
OR2X2 U2190  (.A ( n1297 ) , .B ( n1296 ) , .Y ( n1365 ));
NAND2X2 U2191  (.A ( n1293 ) , .B ( n1292 ) , .Y ( n1295 ));
AOI21X4 U2192  (.A0 ( n1365 ) , .A1 ( n1367 ) , .B0 ( n1298 ) , .Y ( n1454 ));
XOR2X4 U2193  (.A ( n1299 ) , .B ( n1454 ) , .Y ( n1351 ));
INVX2 U2194  (.A ( n1301 ) , .Y ( n1303 ));
NAND2X2 U2195  (.A ( n1707 ) , .B ( n1315 ) , .Y ( n1348 ));
XOR2X1 U2196  (.A ( n1307 ) , .B ( n1348 ) , .Y ( n1309 ));
INVX2 U2197  (.A ( n1308 ) , .Y ( n1311 ));
INVX2 U2198  (.A ( n1309 ) , .Y ( n1310 ));
NAND2X2 U2199  (.A ( n1311 ) , .B ( n1310 ) , .Y ( n1334 ));
NAND2X2 U2200  (.A ( n1312 ) , .B ( n1334 ) , .Y ( n1344 ));
AND2X2 U2201  (.A ( n1582 ) , .B ( n2702 ) , .Y ( n1347 ));
INVX2 U2202  (.A ( n2702 ) , .Y ( n1610 ));
OAI21X1 U2203  (.A0 ( n1610 ) , .A1 ( n1474 ) , .B0 ( n1313 ) , .Y ( n1314 ));
NAND2X2 U2204  (.A ( n1463 ) , .B ( n1314 ) , .Y ( n1320 ));
INVX2 U2205  (.A ( n1707 ) , .Y ( n2698 ));
AND3X2 U2206  (.A ( n1317 ) , .B ( n1316 ) , .C ( n1315 ) , .Y ( n1318 ));
NAND2BX2 U2207  (.AN ( n1320 ) , .B ( n1318 ) , .Y ( n1464 ));
OAI211X2 U2208  (.A0 ( n1321 ) , .A1 ( n1348 ) , .B0 ( n1320 ) , .C0 ( n1319 ) , .Y ( n1322 ));
AOI21X4 U2209  (.A0 ( n1326 ) , .A1 ( n1325 ) , .B0 ( n1324 ) , .Y ( n1328 ));
NAND2X2 U2210  (.A ( n1327 ) , .B ( n1328 ) , .Y ( n1341 ));
INVX2 U2211  (.A ( n1327 ) , .Y ( n1330 ));
NAND2X4 U2212  (.A ( n1330 ) , .B ( n1329 ) , .Y ( n1343 ));
AND2X2 U2213  (.A ( n1341 ) , .B ( n1343 ) , .Y ( n1331 ));
INVX2 U2214  (.A ( n1332 ) , .Y ( n1336 ));
NAND2X4 U2215  (.A ( n1340 ) , .B ( n1339 ) , .Y ( n1361 ));
NAND2X2 U2216  (.A ( n1506 ) , .B ( n1507 ) , .Y ( n1396 ));
NOR2X2 U2217  (.A ( n1367 ) , .B ( n1355 ) , .Y ( n1392 ));
INVX2 U2218  (.A ( n1375 ) , .Y ( n1358 ));
MXI2X1 U2219  (.A ( n1375 ) , .B ( n1356 ) , .S0 ( n1376 ) , .Y ( n1364 ));
OA21X2 U2220  (.A0 ( n1374 ) , .A1 ( n1358 ) , .B0 ( n1357 ) , .Y ( n1363 ));
NAND4X2 U2221  (.A ( n1361 ) , .B ( n1360 ) , .C ( n1359 ) , .D ( n1375 ) , .Y ( n1379 ));
AND2X6 U2222  (.A ( n1392 ) , .B ( n1393 ) , .Y ( n1400 ));
NAND2X2 U2223  (.A ( n1366 ) , .B ( n1365 ) , .Y ( n1368 ));
NAND2BX4 U2224  (.AN ( n1385 ) , .B ( n1383 ) , .Y ( n1409 ));
INVX2 U2225  (.A ( n1383 ) , .Y ( n1384 ));
NAND2X4 U2226  (.A ( n1388 ) , .B ( n1386 ) , .Y ( n1391 ));
INVX2 U2227  (.A ( n1392 ) , .Y ( n1395 ));
XOR2X4 U2228  (.A ( n1396 ) , .B ( n1505 ) , .Y ( n1399 ));
INVX4 U2229  (.A ( n1399 ) , .Y ( n1397 ));
NAND2BX4 U2230  (.AN ( n1398 ) , .B ( n1397 ) , .Y ( n1501 ));
NAND2X2 U2231  (.A ( n1399 ) , .B ( n1398 ) , .Y ( n1483 ));
NAND2X2 U2232  (.A ( n1501 ) , .B ( n1483 ) , .Y ( n1419 ));
INVX4 U2233  (.A ( n1400 ) , .Y ( n1404 ));
XOR2X8 U2234  (.A ( n1402 ) , .B ( n1401 ) , .Y ( n1432 ));
NAND2X4 U2235  (.A ( n1432 ) , .B ( n1433 ) , .Y ( n1437 ));
INVX2 U2236  (.A ( n1407 ) , .Y ( n1408 ));
NAND2X4 U2237  (.A ( n1437 ) , .B ( n1415 ) , .Y ( n1439 ));
INVXL U2238  (.A ( n1412 ) , .Y ( n1413 ));
NAND2X2 U2239  (.A ( n1121 ) , .B ( n1412 ) , .Y ( n1528 ));
AOI2BB2X2 U2240  (.B0 ( n1414 ) , .B1 ( n1413 ) , .A0N ( n1528 ) , .A1N ( n1802 ) , .Y ( n1440 ));
INVX2 U2241  (.A ( n1415 ) , .Y ( n1416 ));
NAND2X4 U2242  (.A ( n1417 ) , .B ( n1416 ) , .Y ( n1438 ));
NAND2X4 U2243  (.A ( n1418 ) , .B ( n1438 ) , .Y ( n1482 ));
XOR2X4 U2244  (.A ( n1419 ) , .B ( n1482 ) , .Y ( n1444 ));
INVX2 U2245  (.A ( n1489 ) , .Y ( n1431 ));
NAND2BX2 U2246  (.AN ( n1431 ) , .B ( n1420 ) , .Y ( n1423 ));
OAI2BB1X1 U2247  (.A0N ( n1427 ) , .A1N ( n1421 ) , .B0 ( n1541 ) , .Y ( n1422 ));
NAND2X2 U2248  (.A ( n1444 ) , .B ( n1445 ) , .Y ( n1906 ));
NAND2XL U2249  (.A ( n1427 ) , .B ( n1820 ) , .Y ( n1428 ));
INVX2 U2250  (.A ( n1432 ) , .Y ( n1435 ));
NAND2X2 U2251  (.A ( n1435 ) , .B ( n1434 ) , .Y ( n1436 ));
AND2X2 U2252  (.A ( n1437 ) , .B ( n1436 ) , .Y ( n2078 ));
NAND3X2 U2253  (.A ( n2078 ) , .B ( n2748 ) , .C ( n1820 ) , .Y ( n1442 ));
XOR2X3 U2254  (.A ( n1441 ) , .B ( n1440 ) , .Y ( n2103 ));
ACHCONX2 U2255  (.A ( n1443 ) , .B ( n1442 ) , .CI ( n2103 ) , .CON ( n1909 ));
NAND2X4 U2256  (.A ( n1906 ) , .B ( n1909 ) , .Y ( n1448 ));
NAND2X2 U2257  (.A ( n1506 ) , .B ( n1555 ) , .Y ( n1452 ));
OAI31X4 U2258  (.A0 ( n1459 ) , .A1 ( n1458 ) , .A2 ( n1056 ) , .B0 ( n1457 ) , .Y ( n1460 ));
OR2X2 U2259  (.A ( n1461 ) , .B ( \intadd_7/SUM[0] ) , .Y ( n1515 ));
NAND2X2 U2260  (.A ( n1461 ) , .B ( \intadd_7/SUM[0] ) , .Y ( n1513 ));
NAND2BX8 U2261  (.AN ( n1468 ) , .B ( n1469 ) , .Y ( n1510 ));
NAND2BX4 U2262  (.AN ( n1469 ) , .B ( n1468 ) , .Y ( n1508 ));
NAND2X2 U2263  (.A ( n1510 ) , .B ( n1508 ) , .Y ( n1470 ));
NAND2X2 U2264  (.A ( n1582 ) , .B ( n1823 ) , .Y ( n1525 ));
INVX2 U2265  (.A ( n1472 ) , .Y ( n1524 ));
OAI21X1 U2266  (.A0 ( n1474 ) , .A1 ( n1049 ) , .B0 ( n1473 ) , .Y ( n1475 ));
OAI21X1 U2267  (.A0 ( n1525 ) , .A1 ( n1524 ) , .B0 ( n1475 ) , .Y ( n1518 ));
NAND2X2 U2268  (.A ( n1528 ) , .B ( n1476 ) , .Y ( n1523 ));
XOR2X1 U2269  (.A ( n1477 ) , .B ( n1522 ) , .Y ( n1480 ));
OR3X2 U2270  (.A ( n1118 ) , .B ( n1487 ) , .C ( n1799 ) , .Y ( n1598 ));
OAI2BB1X1 U2271  (.A0N ( n1598 ) , .A1N ( n1494 ) , .B0 ( n1491 ) , .Y ( n1496 ));
NAND2BX2 U2272  (.AN ( n1118 ) , .B ( n1492 ) , .Y ( n1493 ));
NAND2X2 U2273  (.A ( n1496 ) , .B ( n1599 ) , .Y ( n1540 ));
XOR2X1 U2274  (.A ( n1540 ) , .B ( n1498 ) , .Y ( n1547 ));
NOR2BX8 U2275  (.AN ( n1931 ) , .B ( n1928 ) , .Y ( n1921 ));
NAND2BX2 U2276  (.AN ( n1501 ) , .B ( n1500 ) , .Y ( n1503 ));
AND3X6 U2277  (.A ( n1504 ) , .B ( n1503 ) , .C ( n1502 ) , .Y ( n1606 ));
INVX4 U2278  (.A ( n1505 ) , .Y ( n1512 ));
INVX2 U2279  (.A ( n1507 ) , .Y ( n1511 ));
AOI21X8 U2280  (.A0 ( n1511 ) , .A1 ( n1510 ) , .B0 ( n1509 ) , .Y ( n1562 ));
OAI21X8 U2281  (.A0 ( n1512 ) , .A1 ( n1567 ) , .B0 ( n1562 ) , .Y ( n1571 ));
INVX2 U2282  (.A ( n1513 ) , .Y ( n1514 ));
OR2X2 U2283  (.A ( n1055 ) , .B ( \intadd_7/SUM[1] ) , .Y ( n1517 ));
XOR2X8 U2284  (.A ( n1571 ) , .B ( n1568 ) , .Y ( n1531 ));
AND2X2 U2285  (.A ( n2699 ) , .B ( n1819 ) , .Y ( n1574 ));
INVX2 U2286  (.A ( n1518 ) , .Y ( n1520 ));
NAND2X2 U2287  (.A ( n1522 ) , .B ( n1523 ) , .Y ( n1519 ));
NAND2X2 U2288  (.A ( n1520 ) , .B ( n1519 ) , .Y ( n1521 ));
NAND2X2 U2289  (.A ( n1526 ) , .B ( n2556 ) , .Y ( n1527 ));
MXI2X1 U2290  (.A ( n1527 ) , .B ( n1526 ) , .S0 ( n1580 ) , .Y ( n1577 ));
XOR2X1 U2291  (.A ( n1577 ) , .B ( n1578 ) , .Y ( n1529 ));
NAND2X2 U2292  (.A ( n1605 ) , .B ( n1733 ) , .Y ( n1535 ));
NAND2X2 U2293  (.A ( n1537 ) , .B ( n1536 ) , .Y ( n1538 ));
AND2X2 U2294  (.A ( a[2] ) , .B ( n2556 ) , .Y ( n1593 ));
NAND2X4 U2295  (.A ( n1921 ) , .B ( n1924 ) , .Y ( n1554 ));
NAND2X2 U2296  (.A ( n1924 ) , .B ( n1927 ) , .Y ( n1553 ));
INVX2 U2297  (.A ( n1550 ) , .Y ( n1551 ));
NAND2X2 U2298  (.A ( n1552 ) , .B ( n1551 ) , .Y ( n1923 ));
AND3X6 U2299  (.A ( n1554 ) , .B ( n1553 ) , .C ( n1923 ) , .Y ( n1888 ));
NAND2X8 U2300  (.A ( n1571 ) , .B ( n1570 ) , .Y ( n1693 ));
NAND2BX2 U2301  (.AN ( n1091 ) , .B ( n1823 ) , .Y ( n1685 ));
INVX2 U2302  (.A ( n1574 ) , .Y ( n1632 ));
OAI22X1 U2303  (.A0 ( n1091 ) , .A1 ( n1802 ) , .B0 ( n1575 ) , .B1 ( n1049 ) , .Y ( n1576 ));
OAI21X1 U2304  (.A0 ( n1685 ) , .A1 ( n1632 ) , .B0 ( n1576 ) , .Y ( n1622 ));
NAND2X2 U2305  (.A ( n1582 ) , .B ( n1581 ) , .Y ( n1629 ));
AND2X2 U2306  (.A ( b[3] ) , .B ( n2556 ) , .Y ( n1628 ));
AND2X2 U2307  (.A ( n1629 ) , .B ( n1628 ) , .Y ( n1583 ));
NAND2X2 U2308  (.A ( n1734 ) , .B ( n1736 ) , .Y ( n1589 ));
INVX2 U2309  (.A ( n1666 ) , .Y ( n1604 ));
NAND2BX2 U2310  (.AN ( n1705 ) , .B ( n2732 ) , .Y ( n1716 ));
NAND3XL U2311  (.A ( n1716 ) , .B ( n1818 ) , .C ( n2732 ) , .Y ( n1591 ));
INVX2 U2312  (.A ( n1594 ) , .Y ( n1596 ));
AND2X2 U2313  (.A ( a[3] ) , .B ( n2556 ) , .Y ( n1653 ));
XOR2X1 U2314  (.A ( n1654 ) , .B ( n1600 ) , .Y ( n1647 ));
XOR2X1 U2315  (.A ( n1602 ) , .B ( n1601 ) , .Y ( n1665 ));
INVX2 U2316  (.A ( n1665 ) , .Y ( n1603 ));
INVX4 U2317  (.A ( n1729 ) , .Y ( n1609 ));
NOR2X2 U2318  (.A ( n1610 ) , .B ( n1686 ) , .Y ( n1618 ));
NAND2X2 U2319  (.A ( n1707 ) , .B ( n2734 ) , .Y ( n2755 ));
NAND2BX2 U2320  (.AN ( n2755 ) , .B ( n1618 ) , .Y ( n1613 ));
NAND2X2 U2321  (.A ( n2733 ) , .B ( n2731 ) , .Y ( n2756 ));
NOR2X2 U2322  (.A ( n2754 ) , .B ( n2756 ) , .Y ( n2751 ));
NAND2BX2 U2323  (.AN ( n2752 ) , .B ( n2751 ) , .Y ( n1615 ));
NAND2BX2 U2324  (.AN ( n2755 ) , .B ( n1614 ) , .Y ( n2758 ));
NAND2X2 U2325  (.A ( n1615 ) , .B ( n2758 ) , .Y ( n1617 ));
CLKXOR2X2 U2326  (.A ( \intadd_7/n1  ) , .B ( n1678 ) , .Y ( n1698 ));
XOR2X1 U2327  (.A ( n1699 ) , .B ( n1698 ) , .Y ( n1619 ));
INVX2 U2328  (.A ( n1622 ) , .Y ( n1623 ));
AND2X2 U2329  (.A ( n2734 ) , .B ( n1819 ) , .Y ( n1636 ));
NAND2X2 U2330  (.A ( n1638 ) , .B ( n1637 ) , .Y ( n1639 ));
NAND2X2 U2331  (.A ( n1748 ) , .B ( n1639 ) , .Y ( n1683 ));
NAND2X4 U2332  (.A ( n1641 ) , .B ( n1642 ) , .Y ( n1728 ));
INVX2 U2333  (.A ( n1642 ) , .Y ( n1643 ));
INVX2 U2334  (.A ( n1731 ) , .Y ( n1674 ));
NAND2X2 U2335  (.A ( n1649 ) , .B ( n1648 ) , .Y ( n1651 ));
NAND2X4 U2336  (.A ( n1651 ) , .B ( n1650 ) , .Y ( n1722 ));
NAND2X2 U2337  (.A ( n1707 ) , .B ( n1820 ) , .Y ( n1761 ));
NAND2X2 U2338  (.A ( n1707 ) , .B ( n1657 ) , .Y ( n1712 ));
NAND2BX2 U2339  (.AN ( n1712 ) , .B ( n2733 ) , .Y ( n1715 ));
XOR2X1 U2340  (.A ( n1722 ) , .B ( n1662 ) , .Y ( n1667 ));
INVX2 U2341  (.A ( n1667 ) , .Y ( n1663 ));
AND2X2 U2342  (.A ( n1668 ) , .B ( n1667 ) , .Y ( n1994 ));
OAI21X8 U2343  (.A0 ( n1888 ) , .A1 ( n1889 ) , .B0 ( n1886 ) , .Y ( n2040 ));
NAND3X2 U2344  (.A ( n1671 ) , .B ( n1670 ) , .C ( n1728 ) , .Y ( n1676 ));
NAND2X2 U2345  (.A ( n1693 ) , .B ( n1699 ) , .Y ( n1677 ));
INVX2 U2346  (.A ( n1698 ) , .Y ( n1692 ));
NAND2BX2 U2347  (.AN ( n1678 ) , .B ( \intadd_7/n1  ) , .Y ( n1696 ));
AND2X2 U2348  (.A ( n1696 ) , .B ( n1695 ) , .Y ( n1690 ));
INVX2 U2349  (.A ( n1681 ) , .Y ( n1684 ));
INVX2 U2350  (.A ( n1683 ) , .Y ( n1680 ));
AND2X2 U2351  (.A ( n1751 ) , .B ( b[5] ) , .Y ( n1744 ));
XOR2X1 U2352  (.A ( n1748 ) , .B ( n1744 ) , .Y ( n1689 ));
NOR3X1 U2353  (.A ( n1802 ) , .B ( n1049 ) , .C ( n1686 ) , .Y ( n1687 ));
NAND2X2 U2354  (.A ( n2734 ) , .B ( n1687 ) , .Y ( n1835 ));
NAND3XL U2355  (.A ( n1835 ) , .B ( n1823 ) , .C ( n2734 ) , .Y ( n1688 ));
INVX2 U2356  (.A ( n1730 ) , .Y ( n1702 ));
NAND2BX2 U2357  (.AN ( n1693 ) , .B ( n1692 ) , .Y ( n1701 ));
AOI2BB1X2 U2358  (.A0N ( n1699 ) , .A1N ( n1698 ) , .B0 ( n1697 ) , .Y ( n1700 ));
NAND2X4 U2359  (.A ( n1701 ) , .B ( n1700 ) , .Y ( n1732 ));
NAND2X2 U2360  (.A ( n1702 ) , .B ( n1732 ) , .Y ( n1703 ));
XOR2X8 U2361  (.A ( n1704 ) , .B ( n1703 ) , .Y ( n1770 ));
XOR2X1 U2362  (.A ( n1760 ) , .B ( n1759 ) , .Y ( n1719 ));
INVX2 U2363  (.A ( n1705 ) , .Y ( n1711 ));
OAI21X1 U2364  (.A0 ( n1707 ) , .A1 ( n1706 ) , .B0 ( n2702 ) , .Y ( n1710 ));
NAND2X2 U2365  (.A ( n1707 ) , .B ( n1818 ) , .Y ( n1709 ));
NAND2X2 U2366  (.A ( n2702 ) , .B ( n1820 ) , .Y ( n1708 ));
NAND2X2 U2367  (.A ( n1709 ) , .B ( n1708 ) , .Y ( n1714 ));
NAND2X2 U2368  (.A ( n1763 ) , .B ( n1713 ) , .Y ( n1812 ));
NAND2X2 U2369  (.A ( n1722 ) , .B ( n1721 ) , .Y ( n1723 ));
NAND3X4 U2370  (.A ( n1737 ) , .B ( n1736 ) , .C ( n1735 ) , .Y ( n1738 ));
INVX2 U2371  (.A ( n1744 ) , .Y ( n1749 ));
NAND2X2 U2372  (.A ( n1746 ) , .B ( n1745 ) , .Y ( n1747 ));
NAND2BX2 U2373  (.AN ( n1830 ) , .B ( n1786 ) , .Y ( n1834 ));
NAND2X2 U2374  (.A ( n1781 ) , .B ( n1779 ) , .Y ( n1753 ));
NAND2X2 U2375  (.A ( n1760 ) , .B ( n1759 ) , .Y ( n1757 ));
NAND2X2 U2376  (.A ( n1757 ) , .B ( n1756 ) , .Y ( n1758 ));
XOR2X1 U2377  (.A ( n1793 ) , .B ( a[6] ) , .Y ( n1764 ));
NAND2BX8 U2378  (.AN ( n1767 ) , .B ( n1765 ) , .Y ( n1816 ));
NAND2X2 U2379  (.A ( n1767 ) , .B ( n1766 ) , .Y ( n1768 ));
INVX2 U2380  (.A ( n1770 ) , .Y ( n1773 ));
INVX2 U2381  (.A ( n1771 ) , .Y ( n1772 ));
INVX2 U2382  (.A ( n1779 ) , .Y ( n1780 ));
INVX2 U2383  (.A ( n1782 ) , .Y ( n1783 ));
OAI21X2 U2384  (.A0 ( n1785 ) , .A1 ( n1784 ) , .B0 ( n1783 ) , .Y ( n1832 ));
INVX2 U2385  (.A ( n1788 ) , .Y ( n1789 ));
NAND2BX2 U2386  (.AN ( n1790 ) , .B ( n1789 ) , .Y ( n1836 ));
AND2X2 U2387  (.A ( n1836 ) , .B ( n1805 ) , .Y ( n1791 ));
MXI2X4 U2388  (.A ( n1792 ) , .B ( n1791 ) , .S0 ( n1806 ) , .Y ( n1853 ));
OAI21X1 U2389  (.A0 ( n1794 ) , .A1 ( a[6] ) , .B0 ( n1793 ) , .Y ( n1796 ));
OR2X2 U2390  (.A ( n1799 ) , .B ( n1049 ) , .Y ( n2118 ));
OAI21X4 U2391  (.A0 ( n1811 ) , .A1 ( n1810 ) , .B0 ( n1809 ) , .Y ( n1842 ));
AND2X2 U2392  (.A ( n2118 ) , .B ( n1818 ) , .Y ( n1846 ));
NAND2X2 U2393  (.A ( n1846 ) , .B ( n1823 ) , .Y ( n1867 ));
AND2X2 U2394  (.A ( n1827 ) , .B ( n1826 ) , .Y ( n1845 ));
CLKXOR2X4 U2395  (.A ( n1842 ) , .B ( n1829 ) , .Y ( n1860 ));
NAND4X2 U2396  (.A ( n1836 ) , .B ( n1835 ) , .C ( n1834 ) , .D ( n1833 ) , .Y ( n1857 ));
NOR2X4 U2397  (.A ( n1860 ) , .B ( n1857 ) , .Y ( n1837 ));
INVX2 U2398  (.A ( n1845 ) , .Y ( n1865 ));
NAND2X8 U2399  (.A ( n1851 ) , .B ( n2115 ) , .Y ( n1873 ));
INVX2 U2400  (.A ( n1854 ) , .Y ( n1855 ));
INVX2 U2401  (.A ( n1857 ) , .Y ( n1858 ));
AND3X2 U2402  (.A ( n2112 ) , .B ( n2117 ) , .C ( n2118 ) , .Y ( n1869 ));
AOI21X6 U2403  (.A0 ( n1871 ) , .A1 ( n1900 ) , .B0 ( n1870 ) , .Y ( n1872 ));
CLKNAND2X12 U2404  (.A ( n1873 ) , .B ( n1872 ) , .Y ( n1898 ));
INVXL U2405  (.A ( a[7] ) , .Y ( n1878 ));
NAND3X2 U2406  (.A ( n1884 ) , .B ( n1883 ) , .C ( n2556 ) , .Y ( n2289 ));
OR2X8 U2407  (.A ( n1898 ) , .B ( n1057 ) , .Y ( n2069 ));
INVX12 U2408  (.A ( n2069 ) , .Y ( n1885 ));
INVX18 U2409  (.A ( n1885 ) , .Y ( n2211 ));
INVX4 U2410  (.A ( n1886 ) , .Y ( n1887 ));
INVX2 U2411  (.A ( n1889 ) , .Y ( n1890 ));
INVX2 U2412  (.A ( n1891 ) , .Y ( n2041 ));
NAND2X8 U2413  (.A ( n1894 ) , .B ( n2056 ) , .Y ( n2116 ));
INVX2 U2414  (.A ( n1895 ) , .Y ( n2080 ));
AND2X2 U2415  (.A ( n2080 ) , .B ( n2082 ) , .Y ( n1896 ));
XOR2X3 U2416  (.A ( n2116 ) , .B ( n1896 ) , .Y ( n2070 ));
NAND2BX2 U2417  (.AN ( n2211 ) , .B ( n2070 ) , .Y ( n1904 ));
INVX2 U2418  (.A ( error ) , .Y ( n1897 ));
NAND2X4 U2419  (.A ( n1898 ) , .B ( n1897 ) , .Y ( n1899 ));
CLKBUFX40 U2420  (.A ( n1899 ) , .Y ( n2214 ));
NAND2X2 U2421  (.A ( n2083 ) , .B ( n2081 ) , .Y ( n1901 ));
NAND2BX4 U2422  (.AN ( n2214 ) , .B ( n2079 ) , .Y ( n1903 ));
NAND3X6 U2423  (.A ( n1905 ) , .B ( n1904 ) , .C ( n1903 ) , .Y ( n2372 ));
INVX2 U2424  (.A ( n1951 ) , .Y ( n1919 ));
INVX2 U2425  (.A ( n2017 ) , .Y ( n2210 ));
INVX2 U2426  (.A ( n2078 ) , .Y ( n2075 ));
NOR2X2 U2427  (.A ( n1910 ) , .B ( n2066 ) , .Y ( n2074 ));
AND2X2 U2428  (.A ( n2075 ) , .B ( n2074 ) , .Y ( n2104 ));
NAND2X2 U2429  (.A ( n2103 ) , .B ( n2104 ) , .Y ( n2108 ));
AND2X2 U2430  (.A ( n2017 ) , .B ( n1911 ) , .Y ( n1934 ));
INVX2 U2431  (.A ( n2106 ) , .Y ( n2002 ));
NAND2X2 U2432  (.A ( n1974 ) , .B ( n1912 ) , .Y ( n1978 ));
OA21X4 U2433  (.A0 ( n2214 ) , .A1 ( n1919 ) , .B0 ( n1915 ) , .Y ( n1917 ));
INVXL U2434  (.A ( n1942 ) , .Y ( n1920 ));
AND2X2 U2435  (.A ( \intadd_4/SUM[0] ) , .B ( n1919 ) , .Y ( n1956 ));
INVX2 U2436  (.A ( n1921 ) , .Y ( n1922 ));
NOR2BX4 U2437  (.AN ( n1922 ) , .B ( n1927 ) , .Y ( n1926 ));
NAND2X2 U2438  (.A ( n1924 ) , .B ( n1923 ) , .Y ( n1925 ));
INVX2 U2439  (.A ( n1928 ) , .Y ( n1929 ));
INVX2 U2440  (.A ( n1931 ) , .Y ( n1932 ));
INVX2 U2441  (.A ( n1936 ) , .Y ( n1937 ));
NAND2X2 U2442  (.A ( n1937 ) , .B ( n2007 ) , .Y ( n1939 ));
OAI21X1 U2443  (.A0 ( n2016 ) , .A1 ( n2002 ) , .B0 ( n1978 ) , .Y ( n1938 ));
AOI21X4 U2444  (.A0 ( n1977 ) , .A1 ( n1939 ) , .B0 ( n1938 ) , .Y ( n1940 ));
OA21X4 U2445  (.A0 ( n2214 ) , .A1 ( n1941 ) , .B0 ( n1940 ) , .Y ( n1945 ));
NAND2X8 U2446  (.A ( n1945 ) , .B ( n1944 ) , .Y ( n2152 ));
INVX2 U2447  (.A ( c[12] ) , .Y ( n2523 ));
INVXL U2448  (.A ( n1949 ) , .Y ( n1950 ));
OR2X2 U2449  (.A ( n2211 ) , .B ( n1952 ) , .Y ( n1954 ));
OR2X2 U2450  (.A ( n2214 ) , .B ( \intadd_4/SUM[0] ) , .Y ( n1953 ));
NAND3X8 U2451  (.A ( n1955 ) , .B ( n1954 ) , .C ( n1953 ) , .Y ( n2540 ));
INVX2 U2452  (.A ( c[11] ) , .Y ( n2548 ));
AND2X2 U2453  (.A ( \intadd_4/SUM[1] ) , .B ( n1956 ) , .Y ( n1972 ));
INVXL U2454  (.A ( n1957 ) , .Y ( n1958 ));
NAND2BX2 U2455  (.AN ( n1960 ) , .B ( n1959 ) , .Y ( n1976 ));
INVX2 U2456  (.A ( n1991 ) , .Y ( n1962 ));
AND2X2 U2457  (.A ( n1992 ) , .B ( n1962 ) , .Y ( n1963 ));
OA21X4 U2458  (.A0 ( n2214 ) , .A1 ( n1967 ) , .B0 ( n1966 ) , .Y ( n1968 ));
INVX2 U2459  (.A ( c[13] ) , .Y ( n2537 ));
OA21X4 U2460  (.A0 ( n2214 ) , .A1 ( n1981 ) , .B0 ( n1980 ) , .Y ( n1982 ));
INVXL U2461  (.A ( n1988 ) , .Y ( n1989 ));
AOI22XL U2462  (.A0 ( n1990 ) , .A1 ( n2076 ) , .B0 ( n1989 ) , .B1 ( n2106 ) , .Y ( n2001 ));
NAND2BX2 U2463  (.AN ( n2069 ) , .B ( n2014 ) , .Y ( n2000 ));
AOI21X1 U2464  (.A0 ( n1993 ) , .A1 ( n1992 ) , .B0 ( n1991 ) , .Y ( n1998 ));
XOR2X1 U2465  (.A ( n1998 ) , .B ( n1997 ) , .Y ( n2039 ));
NAND2BX2 U2466  (.AN ( n2214 ) , .B ( n2039 ) , .Y ( n1999 ));
NAND3X6 U2467  (.A ( n2001 ) , .B ( n2000 ) , .C ( n1999 ) , .Y ( n2321 ));
INVX2 U2468  (.A ( c[3] ) , .Y ( n2664 ));
NAND2X2 U2469  (.A ( n2321 ) , .B ( n2664 ) , .Y ( n2035 ));
NAND2BX2 U2470  (.AN ( n2211 ) , .B ( n2213 ) , .Y ( n2223 ));
OAI21XL U2471  (.A0 ( n2290 ) , .A1 ( n2003 ) , .B0 ( n2002 ) , .Y ( n2006 ));
NOR2XL U2472  (.A ( n2290 ) , .B ( n2020 ) , .Y ( n2005 ));
MXI2X1 U2473  (.A ( n2006 ) , .B ( n2005 ) , .S0 ( n2004 ) , .Y ( n2224 ));
NAND2BX2 U2474  (.AN ( n2214 ) , .B ( n2007 ) , .Y ( n2222 ));
NAND4X4 U2475  (.A ( n2223 ) , .B ( n2224 ) , .C ( c[1] ) , .D ( n2222 ) , .Y ( n2027 ));
NAND2BX4 U2476  (.AN ( n2211 ) , .B ( n2007 ) , .Y ( n2031 ));
INVXL U2477  (.A ( n2008 ) , .Y ( n2013 ));
INVXL U2478  (.A ( n2009 ) , .Y ( n2010 ));
NAND3XL U2479  (.A ( n2076 ) , .B ( n2012 ) , .C ( n2011 ) , .Y ( n2029 ));
NAND2XL U2480  (.A ( n2013 ) , .B ( n2106 ) , .Y ( n2028 ));
AND3XL U2481  (.A ( n2029 ) , .B ( c[2] ) , .C ( n2028 ) , .Y ( n2015 ));
NAND2BX4 U2482  (.AN ( n2214 ) , .B ( n2014 ) , .Y ( n2030 ));
NAND3X2 U2483  (.A ( n2031 ) , .B ( n2015 ) , .C ( n2030 ) , .Y ( n2026 ));
OAI22X1 U2484  (.A0 ( n2018 ) , .A1 ( c[1] ) , .B0 ( n2017 ) , .B1 ( c[0] ) , .Y ( n2019 ));
NAND2BX2 U2485  (.AN ( n2211 ) , .B ( n2019 ) , .Y ( n2023 ));
INVXL U2486  (.A ( n2224 ) , .Y ( n2021 ));
NOR2XL U2487  (.A ( n2020 ) , .B ( n2556 ) , .Y ( n2212 ));
INVX2 U2488  (.A ( c[0] ) , .Y ( n2483 ));
AOI22XL U2489  (.A0 ( n2021 ) , .A1 ( n2672 ) , .B0 ( n2212 ) , .B1 ( n2483 ) , .Y ( n2022 ));
OAI2B11X2 U2490  (.A1N ( n2024 ) , .A0 ( n2214 ) , .B0 ( n2023 ) , .C0 ( n2022 ) , .Y ( n2025 ));
NAND3X4 U2491  (.A ( n2027 ) , .B ( n2026 ) , .C ( n2025 ) , .Y ( n2034 ));
NAND2X2 U2492  (.A ( n2337 ) , .B ( n2582 ) , .Y ( n2033 ));
NAND3X4 U2493  (.A ( n2035 ) , .B ( n2034 ) , .C ( n2033 ) , .Y ( n2050 ));
AOI22XL U2494  (.A0 ( n2038 ) , .A1 ( n2051 ) , .B0 ( n2037 ) , .B1 ( n2106 ) , .Y ( n2047 ));
NAND2X2 U2495  (.A ( n2042 ) , .B ( n2041 ) , .Y ( n2043 ));
XOR2X1 U2496  (.A ( n2044 ) , .B ( n2043 ) , .Y ( n2054 ));
NAND2BX2 U2497  (.AN ( n2214 ) , .B ( n2054 ) , .Y ( n2045 ));
NAND3X6 U2498  (.A ( n2047 ) , .B ( n2046 ) , .C ( n2045 ) , .Y ( n2313 ));
NAND2BX2 U2499  (.AN ( n2313 ) , .B ( c[4] ) , .Y ( n2049 ));
NAND2BX2 U2500  (.AN ( n2321 ) , .B ( c[3] ) , .Y ( n2048 ));
NAND3X4 U2501  (.A ( n2050 ) , .B ( n2049 ) , .C ( n2048 ) , .Y ( n2094 ));
INVX2 U2502  (.A ( c[4] ) , .Y ( n2580 ));
AOI22XL U2503  (.A0 ( n2053 ) , .A1 ( n2076 ) , .B0 ( n2052 ) , .B1 ( n2106 ) , .Y ( n2061 ));
AND2X2 U2504  (.A ( n2056 ) , .B ( n2055 ) , .Y ( n2058 ));
XOR2X1 U2505  (.A ( n2058 ) , .B ( n2057 ) , .Y ( n2068 ));
NAND2BX2 U2506  (.AN ( n2214 ) , .B ( n2068 ) , .Y ( n2059 ));
INVX2 U2507  (.A ( c[5] ) , .Y ( n2656 ));
AOI22X2 U2508  (.A0 ( n2580 ) , .A1 ( n2313 ) , .B0 ( n2329 ) , .B1 ( n2656 ) , .Y ( n2093 ));
INVX2 U2509  (.A ( n2062 ) , .Y ( n2065 ));
AOI22XL U2510  (.A0 ( n2067 ) , .A1 ( n2066 ) , .B0 ( n2106 ) , .B1 ( n2065 ) , .Y ( n2073 ));
NAND2BX2 U2511  (.AN ( n2069 ) , .B ( n2068 ) , .Y ( n2072 ));
NAND2BX2 U2512  (.AN ( n2214 ) , .B ( n2070 ) , .Y ( n2071 ));
NAND2BX2 U2513  (.AN ( n2382 ) , .B ( c[6] ) , .Y ( n2091 ));
NAND2BX2 U2514  (.AN ( n2329 ) , .B ( c[5] ) , .Y ( n2090 ));
XOR2X1 U2515  (.A ( n2075 ) , .B ( n2074 ) , .Y ( n2077 ));
NAND2X2 U2516  (.A ( n2077 ) , .B ( n2076 ) , .Y ( n2097 ));
NAND2BX4 U2517  (.AN ( n2211 ) , .B ( n2079 ) , .Y ( n2100 ));
AND2X2 U2518  (.A ( n2081 ) , .B ( n2080 ) , .Y ( n2085 ));
NAND2X2 U2519  (.A ( n2086 ) , .B ( n2112 ) , .Y ( n2087 ));
XOR2X4 U2520  (.A ( n2088 ) , .B ( n2087 ) , .Y ( n2102 ));
NAND3X4 U2521  (.A ( n2089 ) , .B ( n2100 ) , .C ( n2098 ) , .Y ( n2127 ));
NAND2BX8 U2522  (.AN ( n2372 ) , .B ( c[7] ) , .Y ( n2101 ));
NAND4X4 U2523  (.A ( n2091 ) , .B ( n2090 ) , .C ( n2127 ) , .D ( n2101 ) , .Y ( n2092 ));
AND3X2 U2524  (.A ( n2100 ) , .B ( n2099 ) , .C ( n2098 ) , .Y ( n2300 ));
NAND2BX2 U2525  (.AN ( n2211 ) , .B ( n2102 ) , .Y ( n2126 ));
INVXL U2526  (.A ( n2118 ) , .Y ( n2119 ));
NAND2BX2 U2527  (.AN ( n2214 ) , .B ( n2123 ) , .Y ( n2124 ));
NAND3X4 U2528  (.A ( n2127 ) , .B ( n2372 ) , .C ( n2503 ) , .Y ( n2128 ));
OA21X4 U2529  (.A0 ( c[9] ) , .A1 ( n2187 ) , .B0 ( n2128 ) , .Y ( n2129 ));
OAI2B11X4 U2530  (.A1N ( n2131 ) , .A0 ( n2300 ) , .B0 ( n2130 ) , .C0 ( n2129 ) , .Y ( n2133 ));
INVX2 U2531  (.A ( c[10] ) , .Y ( n2632 ));
OAI22X4 U2532  (.A0 ( n2540 ) , .A1 ( n2548 ) , .B0 ( n2445 ) , .B1 ( n2632 ) , .Y ( n2137 ));
INVX2 U2533  (.A ( n2135 ) , .Y ( n2136 ));
NAND3X2 U2534  (.A ( n2140 ) , .B ( n2139 ) , .C ( n2138 ) , .Y ( n2141 ));
OAI2BB1X4 U2535  (.A0N ( n2146 ) , .A1N ( n2145 ) , .B0 ( n2144 ) , .Y ( n2161 ));
MXI2X1 U2536  (.A ( c[6] ) , .B ( n2382 ) , .S0 ( n2218 ) , .Y ( n2237 ));
NAND2X2 U2537  (.A ( n2505 ) , .B ( n2632 ) , .Y ( n2147 ));
INVX4 U2538  (.A ( n2277 ) , .Y ( n2241 ));
MXI2X2 U2539  (.A ( n2523 ) , .B ( n2522 ) , .S0 ( n2189 ) , .Y ( n2148 ));
INVXL U2540  (.A ( n2149 ) , .Y ( n2150 ));
NOR2X2 U2541  (.A ( n2153 ) , .B ( n2152 ) , .Y ( n2154 ));
NAND3X6 U2542  (.A ( n2172 ) , .B ( n2601 ) , .C ( n2156 ) , .Y ( n2179 ));
MXI2X2 U2543  (.A ( n2158 ) , .B ( n2157 ) , .S0 ( n2189 ) , .Y ( n2159 ));
INVX2 U2544  (.A ( n2540 ) , .Y ( n2519 ));
XOR2X8 U2545  (.A ( n2164 ) , .B ( n2175 ) , .Y ( n2203 ));
OA22X2 U2546  (.A0 ( n2219 ) , .A1 ( n2269 ) , .B0 ( n2259 ) , .B1 ( n2208 ) , .Y ( n2192 ));
NAND2X4 U2547  (.A ( n2172 ) , .B ( n2171 ) , .Y ( n2173 ));
NAND3X4 U2548  (.A ( n2183 ) , .B ( n2549 ) , .C ( n2173 ) , .Y ( n2197 ));
INVX2 U2549  (.A ( n2175 ) , .Y ( n2176 ));
AND2X2 U2550  (.A ( n2182 ) , .B ( n2181 ) , .Y ( n2185 ));
NOR2X2 U2551  (.A ( n2171 ) , .B ( n2185 ) , .Y ( n2186 ));
INVXL U2552  (.A ( c[9] ) , .Y ( n2188 ));
MXI2X1 U2553  (.A ( n2188 ) , .B ( n2187 ) , .S0 ( n2189 ) , .Y ( n2232 ));
MXI2X1 U2554  (.A ( n2131 ) , .B ( n2300 ) , .S0 ( n2189 ) , .Y ( n2244 ));
INVX2 U2555  (.A ( n2229 ) , .Y ( n2190 ));
NAND2X2 U2556  (.A ( n2278 ) , .B ( n2190 ) , .Y ( n2191 ));
MXI2X1 U2557  (.A ( c[2] ) , .B ( n2337 ) , .S0 ( n2218 ) , .Y ( n2248 ));
NOR2X2 U2558  (.A ( n2259 ) , .B ( n2209 ) , .Y ( n2194 ));
OA22X2 U2559  (.A0 ( n2208 ) , .A1 ( n2269 ) , .B0 ( n2247 ) , .B1 ( n2204 ) , .Y ( n2205 ));
OA22X2 U2560  (.A0 ( n2209 ) , .A1 ( n2269 ) , .B0 ( n2239 ) , .B1 ( n2208 ) , .Y ( n2228 ));
INVXL U2561  (.A ( n2212 ) , .Y ( n2216 ));
OA22X2 U2562  (.A0 ( n2220 ) , .A1 ( n2439 ) , .B0 ( n2247 ) , .B1 ( n2219 ) , .Y ( n2227 ));
AND2X2 U2563  (.A ( n2221 ) , .B ( n2277 ) , .Y ( n2249 ));
NAND3X2 U2564  (.A ( n2249 ) , .B ( n2275 ) , .C ( n2236 ) , .Y ( n2225 ));
AND3X2 U2565  (.A ( n2251 ) , .B ( n2252 ) , .C ( n2225 ) , .Y ( n2226 ));
MXI2X1 U2566  (.A ( n2238 ) , .B ( n2237 ) , .S0 ( n2277 ) , .Y ( n2265 ));
OA22X2 U2567  (.A0 ( n2240 ) , .A1 ( n2439 ) , .B0 ( n2239 ) , .B1 ( n2265 ) , .Y ( n2255 ));
OA22X2 U2568  (.A0 ( n2258 ) , .A1 ( n2269 ) , .B0 ( n2268 ) , .B1 ( n2247 ) , .Y ( n2254 ));
NAND3X2 U2569  (.A ( n2275 ) , .B ( n2249 ) , .C ( n2248 ) , .Y ( n2250 ));
AND3X2 U2570  (.A ( n2252 ) , .B ( n2251 ) , .C ( n2250 ) , .Y ( n2253 ));
NAND3X4 U2571  (.A ( n2255 ) , .B ( n2254 ) , .C ( n2253 ) , .Y ( n2256 ));
NAND2BX2 U2572  (.AN ( n2259 ) , .B ( n2258 ) , .Y ( n2263 ));
NAND2X4 U2573  (.A ( n2264 ) , .B ( n2411 ) , .Y ( n2317 ));
INVX2 U2574  (.A ( n2265 ) , .Y ( n2272 ));
NAND2BX2 U2575  (.AN ( n2269 ) , .B ( n2268 ) , .Y ( n2270 ));
OAI211X2 U2576  (.A0 ( n2259 ) , .A1 ( n2272 ) , .B0 ( n2271 ) , .C0 ( n2270 ) , .Y ( n2273 ));
NAND2X8 U2577  (.A ( n2325 ) , .B ( n2324 ) , .Y ( n2374 ));
NAND2X2 U2578  (.A ( n2278 ) , .B ( n2277 ) , .Y ( n2282 ));
AND3X2 U2579  (.A ( n2282 ) , .B ( n2281 ) , .C ( n2247 ) , .Y ( n2285 ));
NAND2X8 U2580  (.A ( n2287 ) , .B ( n2297 ) , .Y ( n2413 ));
NAND2X2 U2581  (.A ( n2690 ) , .B ( n2293 ) , .Y ( n2742 ));
MXI2X1 U2582  (.A ( c[8] ) , .B ( n2301 ) , .S0 ( n2621 ) , .Y ( n2302 ));
NAND2X4 U2583  (.A ( n2320 ) , .B ( n2306 ) , .Y ( n2312 ));
OAI21X2 U2584  (.A0 ( n2307 ) , .A1 ( n2550 ) , .B0 ( n2296 ) , .Y ( n2309 ));
NAND2X4 U2585  (.A ( n2309 ) , .B ( n2308 ) , .Y ( n2311 ));
MXI2X1 U2586  (.A ( n2580 ) , .B ( n2314 ) , .S0 ( n2621 ) , .Y ( n2364 ));
INVX2 U2587  (.A ( n2317 ) , .Y ( n2315 ));
OAI21X2 U2588  (.A0 ( n2316 ) , .A1 ( n2332 ) , .B0 ( n2315 ) , .Y ( n2319 ));
OAI22X1 U2589  (.A0 ( n2317 ) , .A1 ( n2296 ) , .B0 ( n2556 ) , .B1 ( n2664 ) , .Y ( n2318 ));
MXI2X1 U2590  (.A ( c[3] ) , .B ( n2321 ) , .S0 ( n2621 ) , .Y ( n2355 ));
INVX2 U2591  (.A ( n2355 ) , .Y ( n2322 ));
INVX2 U2592  (.A ( n2296 ) , .Y ( n2564 ));
NOR2BX1 U2593  (.AN ( c[5] ) , .B ( n2556 ) , .Y ( n2326 ));
MXI2X1 U2594  (.A ( n2656 ) , .B ( n2330 ) , .S0 ( n2621 ) , .Y ( n2359 ));
MXI2X1 U2595  (.A ( c[2] ) , .B ( n2337 ) , .S0 ( n2621 ) , .Y ( n2351 ));
INVX2 U2596  (.A ( n2338 ) , .Y ( n2344 ));
INVX2 U2597  (.A ( n2340 ) , .Y ( n2341 ));
AND2X2 U2598  (.A ( n2345 ) , .B ( n2341 ) , .Y ( n2343 ));
AOI22X2 U2599  (.A0 ( n2341 ) , .A1 ( n2564 ) , .B0 ( c[1] ) , .B1 ( n2692 ) , .Y ( n2342 ));
OAI21X6 U2600  (.A0 ( n2344 ) , .A1 ( n2343 ) , .B0 ( n2342 ) , .Y ( n2481 ));
MXI2X1 U2601  (.A ( c[1] ) , .B ( n2348 ) , .S0 ( n2621 ) , .Y ( n2349 ));
NAND2X4 U2602  (.A ( n2350 ) , .B ( n2480 ) , .Y ( n2493 ));
INVX2 U2603  (.A ( n2351 ) , .Y ( n2352 ));
NAND2X2 U2604  (.A ( n2353 ) , .B ( n2352 ) , .Y ( n2491 ));
NAND2X2 U2605  (.A ( n2356 ) , .B ( n2355 ) , .Y ( n2484 ));
NAND2X8 U2606  (.A ( n2486 ) , .B ( n2484 ) , .Y ( n2426 ));
INVX2 U2607  (.A ( n2358 ) , .Y ( n2360 ));
INVX2 U2608  (.A ( n2363 ) , .Y ( n2366 ));
INVX2 U2609  (.A ( n2364 ) , .Y ( n2365 ));
NAND2X4 U2610  (.A ( n2366 ) , .B ( n2365 ) , .Y ( n2456 ));
NAND2X4 U2611  (.A ( n2403 ) , .B ( n2428 ) , .Y ( n2383 ));
NAND2X2 U2612  (.A ( n2367 ) , .B ( n2368 ) , .Y ( n2370 ));
OR2X2 U2613  (.A ( n2371 ) , .B ( n2296 ) , .Y ( n2389 ));
AND3X2 U2614  (.A ( n2389 ) , .B ( n2395 ) , .C ( n2390 ) , .Y ( n2373 ));
NAND2X4 U2615  (.A ( n2375 ) , .B ( n2376 ) , .Y ( n2381 ));
AND3X6 U2616  (.A ( n2381 ) , .B ( n2380 ) , .C ( n2379 ) , .Y ( n2385 ));
NAND4X6 U2617  (.A ( n2384 ) , .B ( n2383 ) , .C ( n2407 ) , .D ( n2423 ) , .Y ( n2399 ));
INVX2 U2618  (.A ( n2386 ) , .Y ( n2387 ));
NAND2BX4 U2619  (.AN ( n2422 ) , .B ( n2407 ) , .Y ( n2398 ));
NOR2X2 U2620  (.A ( n2392 ) , .B ( n2391 ) , .Y ( n2393 ));
NAND2X2 U2621  (.A ( n2394 ) , .B ( n2393 ) , .Y ( n2397 ));
INVX2 U2622  (.A ( n2395 ) , .Y ( n2396 ));
NAND2X4 U2623  (.A ( n2401 ) , .B ( n2426 ) , .Y ( n2402 ));
NAND2BX2 U2624  (.AN ( n2403 ) , .B ( n2402 ) , .Y ( n2404 ));
AND2X2 U2625  (.A ( n2407 ) , .B ( n2406 ) , .Y ( n2408 ));
AND2X4 U2626  (.A ( n2694 ) , .B ( n2677 ) , .Y ( n2454 ));
NAND2BX8 U2627  (.AN ( n2413 ) , .B ( n2415 ) , .Y ( n2444 ));
AOI2BB2X2 U2628  (.B0 ( c[9] ) , .B1 ( n2692 ) , .A0N ( n2415 ) , .A1N ( n2296 ) , .Y ( n2416 ));
INVX2 U2629  (.A ( n2420 ) , .Y ( n2419 ));
NAND2X2 U2630  (.A ( n2423 ) , .B ( n2422 ) , .Y ( n2424 ));
XOR2X4 U2631  (.A ( n2425 ) , .B ( n2424 ) , .Y ( n2673 ));
CLKXOR2X4 U2632  (.A ( n2431 ) , .B ( n2430 ) , .Y ( n2654 ));
NAND2X8 U2633  (.A ( n2436 ) , .B ( n2435 ) , .Y ( n2464 ));
INVXL U2634  (.A ( n2461 ) , .Y ( n2446 ));
NAND3X2 U2635  (.A ( n2462 ) , .B ( n2448 ) , .C ( n2447 ) , .Y ( n2449 ));
XOR2X8 U2636  (.A ( n2450 ) , .B ( n2449 ) , .Y ( n2588 ));
NAND3X8 U2637  (.A ( n2454 ) , .B ( n2451 ) , .C ( n2588 ) , .Y ( n2680 ));
NAND3X4 U2638  (.A ( n2588 ) , .B ( n2591 ) , .C ( n2453 ) , .Y ( n2488 ));
CLKNAND2X12 U2639  (.A ( n2588 ) , .B ( n2688 ) , .Y ( n2678 ));
NAND3X8 U2640  (.A ( n2680 ) , .B ( n2488 ) , .C ( n2678 ) , .Y ( n2510 ));
AND2X2 U2641  (.A ( n2456 ) , .B ( n2455 ) , .Y ( n2457 ));
INVX2 U2642  (.A ( n2683 ) , .Y ( n2647 ));
NAND3X8 U2643  (.A ( n2625 ) , .B ( n2686 ) , .C ( n2674 ) , .Y ( n2642 ));
NAND2X2 U2644  (.A ( n2469 ) , .B ( n2468 ) , .Y ( n2470 ));
CLKXOR2X2 U2645  (.A ( n2482 ) , .B ( n2481 ) , .Y ( n2657 ));
CLKXOR2X2 U2646  (.A ( n2487 ) , .B ( n2486 ) , .Y ( n2679 ));
AOI22X2 U2647  (.A0 ( n2490 ) , .A1 ( n2683 ) , .B0 ( n2489 ) , .B1 ( n2654 ) , .Y ( n2498 ));
INVX2 U2648  (.A ( n2680 ) , .Y ( n2496 ));
CLKXOR2X2 U2649  (.A ( n2495 ) , .B ( n2494 ) , .Y ( n2636 ));
INVX2 U2650  (.A ( n2677 ) , .Y ( n2638 ));
NAND3X4 U2651  (.A ( n2680 ) , .B ( n2686 ) , .C ( n2633 ) , .Y ( n2600 ));
NOR2X2 U2652  (.A ( n2568 ) , .B ( n2550 ) , .Y ( n2517 ));
BUFX2 U2653  (.A ( n2504 ) , .Y ( n2595 ));
NAND3X2 U2654  (.A ( n2601 ) , .B ( n2595 ) , .C ( n2627 ) , .Y ( n2561 ));
NAND3XL U2655  (.A ( n2597 ) , .B ( n2549 ) , .C ( n2628 ) , .Y ( n2507 ));
NAND3X2 U2656  (.A ( n2508 ) , .B ( n2673 ) , .C ( n2683 ) , .Y ( n2509 ));
NAND2X8 U2657  (.A ( n2510 ) , .B ( n2627 ) , .Y ( n2623 ));
AOI21X8 U2658  (.A0 ( n2513 ) , .A1 ( n2512 ) , .B0 ( n2511 ) , .Y ( n2603 ));
AOI22X4 U2659  (.A0 ( n2603 ) , .A1 ( n2598 ) , .B0 ( n2642 ) , .B1 ( n2600 ) , .Y ( n2736 ));
NOR2X6 U2660  (.A ( n2521 ) , .B ( n2556 ) , .Y ( n2617 ));
NOR2X2 U2661  (.A ( n2530 ) , .B ( n2529 ) , .Y ( n2553 ));
NOR3X2 U2662  (.A ( n2570 ) , .B ( n2549 ) , .C ( n2571 ) , .Y ( n2738 ));
NOR2X2 U2663  (.A ( n2554 ) , .B ( c[14] ) , .Y ( n2567 ));
NOR2X2 U2664  (.A ( n2550 ) , .B ( n2655 ) , .Y ( n2599 ));
AOI21X1 U2665  (.A0 ( n2617 ) , .A1 ( n2610 ) , .B0 ( n2614 ) , .Y ( n2560 ));
NOR2BXL U2666  (.AN ( c[14] ) , .B ( n2556 ) , .Y ( n2557 ));
OR2X2 U2667  (.A ( n2558 ) , .B ( n2557 ) , .Y ( n2613 ));
NAND3XL U2668  (.A ( n2568 ) , .B ( n2567 ) , .C ( n2599 ) , .Y ( n2569 ));
MXI2X2 U2669  (.A ( n2573 ) , .B ( n2572 ) , .S0 ( n2736 ) , .Y ( n2574 ));
OAI22X1 U2670  (.A0 ( n2673 ) , .A1 ( n2675 ) , .B0 ( n2674 ) , .B1 ( n2677 ) , .Y ( n2587 ));
OAI21X1 U2671  (.A0 ( n2684 ) , .A1 ( n2583 ) , .B0 ( n2654 ) , .Y ( n2586 ));
OAI22X4 U2672  (.A0 ( n2695 ) , .A1 ( n2591 ) , .B0 ( n2590 ) , .B1 ( n2692 ) , .Y ( n2746 ));
NOR2XL U2673  (.A ( n2608 ) , .B ( n2609 ) , .Y ( mac_out[13] ));
INVXL U2674  (.A ( n2611 ) , .Y ( n2612 ));
AO21X2 U2675  (.A0 ( n2617 ) , .A1 ( n2616 ) , .B0 ( n2615 ) , .Y ( n2618 ));
OAI22X2 U2676  (.A0 ( n2647 ) , .A1 ( n2674 ) , .B0 ( n2675 ) , .B1 ( n2679 ) , .Y ( n2635 ));
OAI22X1 U2677  (.A0 ( n2680 ) , .A1 ( n2657 ) , .B0 ( n2678 ) , .B1 ( n2676 ) , .Y ( n2634 ));
AOI211X4 U2678  (.A0 ( n2684 ) , .A1 ( n2636 ) , .B0 ( n2635 ) , .C0 ( n2634 ) , .Y ( n2637 ));
MXI2X1 U2679  (.A ( n2719 ) , .B ( n2672 ) , .S0 ( n2655 ) , .Y ( n1010 ));
OAI22X1 U2680  (.A0 ( n2676 ) , .A1 ( n2675 ) , .B0 ( n2674 ) , .B1 ( n2673 ) , .Y ( n2682 ));
AOI211X4 U2681  (.A0 ( n2684 ) , .A1 ( n2683 ) , .B0 ( n2682 ) , .C0 ( n2681 ) , .Y ( n2685 ));
AOI22X2 U2682  (.A0 ( n2691 ) , .A1 ( n2690 ) , .B0 ( n2689 ) , .B1 ( n2688 ) , .Y ( n2693 ));
OAI22X4 U2683  (.A0 ( n2695 ) , .A1 ( n2694 ) , .B0 ( n2693 ) , .B1 ( n2692 ) , .Y ( n2747 ));
AOI2BB1X2 U2684  (.A0N ( n2697 ) , .A1N ( n2706 ) , .B0 ( n2696 ) , .Y ( n2705 ));
AOI21X1 U2685  (.A0 ( n2705 ) , .A1 ( n2704 ) , .B0 ( n2710 ) , .Y ( \intadd_7/B[0] ));
XOR2X1 U2686  (.A ( n2710 ) , .B ( n2709 ) , .Y ( \intadd_7/A[1] ));
NOR2XL U2687  (.A ( n2608 ) , .B ( n2711 ) , .Y ( mac_out[3] ));
NOR2XL U2688  (.A ( n2608 ) , .B ( n2712 ) , .Y ( mac_out[2] ));
NOR2XL U2689  (.A ( n2608 ) , .B ( n2713 ) , .Y ( mac_out[11] ));
NOR2XL U2690  (.A ( n2608 ) , .B ( n2714 ) , .Y ( mac_out[10] ));
NOR2XL U2691  (.A ( n2608 ) , .B ( n2715 ) , .Y ( mac_out[7] ));
NOR2XL U2692  (.A ( n2608 ) , .B ( n2716 ) , .Y ( mac_out[6] ));
NOR2XL U2693  (.A ( n2608 ) , .B ( n2717 ) , .Y ( mac_out[5] ));
NOR2XL U2694  (.A ( n2608 ) , .B ( n2718 ) , .Y ( mac_out[4] ));
NOR2XL U2695  (.A ( n2608 ) , .B ( n2719 ) , .Y ( mac_out[1] ));
NOR2XL U2696  (.A ( n2608 ) , .B ( n2720 ) , .Y ( mac_out[0] ));
NOR2BXL U2697  (.AN ( clk ) , .B ( clk ) , .Y ( n2721 ));
MX2XL U2698  (.A ( n2556 ) , .B ( clk ) , .S0 ( n2721 ) , .Y ( n1028 ));
MX2XL U2699  (.A ( a[14] ) , .B ( in_a[14] ) , .S0 ( n2749 ) , .Y ( n1026 ));
NOR2XL U2700  (.A ( n2742 ) , .B ( n2722 ) , .Y ( n2723 ));
NOR4XL U2701  (.A ( n2726 ) , .B ( n2725 ) , .C ( n2724 ) , .D ( n2723 ) , .Y ( n2727 ));
NOR2XL U2702  (.A ( n2608 ) , .B ( n2727 ) , .Y ( mac_out[12] ));
AOI21XL U2703  (.A0 ( n2729 ) , .A1 ( c[15] ) , .B0 ( n2728 ) , .Y ( n2730 ));
NOR2XL U2704  (.A ( n2608 ) , .B ( n2730 ) , .Y ( mac_out[15] ));
AOI22XL U2705  (.A0 ( n2734 ) , .A1 ( n2733 ) , .B0 ( n2732 ) , .B1 ( n2731 ) , .Y ( n2735 ));
INVXL U2706  (.A ( n2736 ) , .Y ( n2737 ));
NAND2XL U2707  (.A ( n2738 ) , .B ( n2737 ) , .Y ( n2739 ));
XOR2XL U2708  (.A ( n2740 ) , .B ( n2739 ) , .Y ( n2743 ));
OAI21XL U2709  (.A0 ( n2743 ) , .A1 ( n2742 ) , .B0 ( n2741 ) , .Y ( n2744 ));
AOI2BB1XL U2710  (.A0N ( n2745 ) , .A1N ( n2744 ) , .B0 ( n2608 ) , .Y ( mac_out[14] ));
NOR2BXL U2711  (.AN ( n2746 ) , .B ( n2608 ) , .Y ( mac_out[9] ));
NOR2BXL U2712  (.AN ( n2747 ) , .B ( n2608 ) , .Y ( mac_out[8] ));
MX2XL U2713  (.A ( a[13] ) , .B ( in_a[13] ) , .S0 ( n1048 ) , .Y ( n1025 ));
MX2XL U2714  (.A ( a[12] ) , .B ( in_a[12] ) , .S0 ( n1048 ) , .Y ( n1024 ));
MX2XL U2715  (.A ( a[11] ) , .B ( in_a[11] ) , .S0 ( n1048 ) , .Y ( n1023 ));
MX2XL U2716  (.A ( b[14] ) , .B ( in_b[14] ) , .S0 ( n1048 ) , .Y ( n1043 ));
MX2XL U2717  (.A ( b[13] ) , .B ( in_b[13] ) , .S0 ( n1048 ) , .Y ( n1042 ));
MX2XL U2718  (.A ( b[12] ) , .B ( in_b[12] ) , .S0 ( n1048 ) , .Y ( n1041 ));
MX2XL U2719  (.A ( b[11] ) , .B ( in_b[11] ) , .S0 ( n1048 ) , .Y ( n1040 ));
MX2XL U2720  (.A ( b[10] ) , .B ( in_b[10] ) , .S0 ( n1048 ) , .Y ( n1039 ));
MX2XL U2721  (.A ( a[10] ) , .B ( in_a[10] ) , .S0 ( n1048 ) , .Y ( n1022 ));
MX2XL U2722  (.A ( n2748 ) , .B ( in_a[0] ) , .S0 ( n1048 ) , .Y ( n1012 ));
MX2XL U2723  (.A ( a[1] ) , .B ( in_a[1] ) , .S0 ( n1048 ) , .Y ( n1013 ));
MX2XL U2724  (.A ( a[2] ) , .B ( in_a[2] ) , .S0 ( n1048 ) , .Y ( n1014 ));
MX2XL U2725  (.A ( a[3] ) , .B ( in_a[3] ) , .S0 ( n1048 ) , .Y ( n1015 ));
MX2XL U2726  (.A ( a[4] ) , .B ( in_a[4] ) , .S0 ( n1048 ) , .Y ( n1016 ));
MX2XL U2727  (.A ( a[5] ) , .B ( in_a[5] ) , .S0 ( n1048 ) , .Y ( n1017 ));
MX2XL U2728  (.A ( a[6] ) , .B ( in_a[6] ) , .S0 ( n1048 ) , .Y ( n1018 ));
MX2XL U2729  (.A ( a[7] ) , .B ( in_a[7] ) , .S0 ( n1048 ) , .Y ( n1019 ));
MX2XL U2730  (.A ( a[8] ) , .B ( in_a[8] ) , .S0 ( n1048 ) , .Y ( n1020 ));
MX2XL U2731  (.A ( a[9] ) , .B ( in_a[9] ) , .S0 ( n1048 ) , .Y ( n1021 ));
MX2XL U2732  (.A ( a[15] ) , .B ( in_a[15] ) , .S0 ( n1048 ) , .Y ( n1027 ));
MX2XL U2733  (.A ( n2750 ) , .B ( in_b[0] ) , .S0 ( n1048 ) , .Y ( n1029 ));
MX2XL U2734  (.A ( b[2] ) , .B ( in_b[2] ) , .S0 ( n1048 ) , .Y ( n1031 ));
MX2XL U2735  (.A ( b[3] ) , .B ( in_b[3] ) , .S0 ( n1048 ) , .Y ( n1032 ));
MX2XL U2736  (.A ( b[4] ) , .B ( in_b[4] ) , .S0 ( n1048 ) , .Y ( n1033 ));
MX2XL U2737  (.A ( b[5] ) , .B ( in_b[5] ) , .S0 ( n1048 ) , .Y ( n1034 ));
MX2XL U2738  (.A ( b[6] ) , .B ( in_b[6] ) , .S0 ( n1048 ) , .Y ( n1035 ));
MX2XL U2739  (.A ( b[8] ) , .B ( in_b[8] ) , .S0 ( n1048 ) , .Y ( n1037 ));
MX2XL U2740  (.A ( b[9] ) , .B ( in_b[9] ) , .S0 ( n1048 ) , .Y ( n1038 ));
MX2XL U2741  (.A ( b[15] ) , .B ( in_b[15] ) , .S0 ( n1048 ) , .Y ( n1044 ));
NAND2BX2 U2742  (.AN ( n2751 ) , .B ( n2758 ) , .Y ( n2753 ));
XNOR2X1 U2743  (.A ( n2753 ) , .B ( n2752 ) , .Y ( \intadd_7/A[2] ));
OAI21X1 U2744  (.A0 ( n2757 ) , .A1 ( n2756 ) , .B0 ( n2755 ) , .Y ( n2759 ));
AND2X2 U2745  (.A ( n2759 ) , .B ( n2758 ) , .Y ( \intadd_7/B[1] ));
endmodule
