module s1238_bench (G3 , G2 , G1 , G0 , blif_reset_net , blif_clk_net , 
    G11 , G10 , G9 , G8 , G7 , G6 , G5 , G4 , G546 , G542 , G552 , 
    G551 , G550 , G549 , G13 , G12 , G539 , G45 , G537 , G535 , 
    G532 , G530 , G548 , G547 );
input  G3 ;
input  G2 ;
input  G1 ;
input  G0 ;
input  blif_reset_net ;
input  blif_clk_net ;
input  G11 ;
input  G10 ;
input  G9 ;
input  G8 ;
input  G7 ;
input  G6 ;
input  G5 ;
input  G4 ;
output G546 ;
output G542 ;
output G552 ;
output G551 ;
output G550 ;
output G549 ;
input  G13 ;
input  G12 ;
output G539 ;
output G45 ;
output G537 ;
output G535 ;
output G532 ;
output G530 ;
output G548 ;
output G547 ;



INV_X0P5B_A9TL40 U98 (.A ( n646 ) , .Y ( n668 ) ) ;
INV_X0P8M_A9TL40 U97 (.A ( n668 ) , .Y ( n667 ) ) ;
INV_X0P5B_A9TL40 U96 (.A ( G11 ) , .Y ( n666 ) ) ;
INV_X1M_A9TL40 U95 (.A ( n666 ) , .Y ( n665 ) ) ;
INV_X0P5B_A9TL40 U94 (.A ( n645 ) , .Y ( n664 ) ) ;
INV_X0P6M_A9TL40 U93 (.A ( n664 ) , .Y ( n663 ) ) ;
INV_X0P5B_A9TL40 U92 (.A ( n643 ) , .Y ( n662 ) ) ;
INV_X0P6M_A9TL40 U91 (.A ( n662 ) , .Y ( n661 ) ) ;
INV_X0P5B_A9TL40 U90 (.A ( n641 ) , .Y ( n660 ) ) ;
INV_X1B_A9TL40 U89 (.A ( n660 ) , .Y ( n659 ) ) ;
INV_X0P5B_A9TL40 U88 (.A ( n639 ) , .Y ( n658 ) ) ;
INV_X0P8M_A9TL40 U87 (.A ( n658 ) , .Y ( n657 ) ) ;
BUF_X1P2M_A9TL40 U86 (.A ( n638 ) , .Y ( n656 ) ) ;
INV_X0P5B_A9TL40 U85 (.A ( n636 ) , .Y ( n655 ) ) ;
INV_X0P7B_A9TL40 U84 (.A ( n655 ) , .Y ( n654 ) ) ;
INV_X0P5B_A9TL40 U83 (.A ( n634 ) , .Y ( n653 ) ) ;
INV_X0P7B_A9TL40 U82 (.Y ( n652 ) , .A ( n653 ) ) ;
INV_X0P5B_A9TL40 U81 (.A ( n632 ) , .Y ( n651 ) ) ;
INV_X0P7B_A9TL40 U80 (.A ( n651 ) , .Y ( n650 ) ) ;
INV_X0P5B_A9TL40 U79 (.A ( n630 ) , .Y ( n649 ) ) ;
INV_X0P8M_A9TL40 U78 (.A ( n649 ) , .Y ( n648 ) ) ;
INV_X0P5B_A9TL40 U77 (.A ( G12 ) , .Y ( n647 ) ) ;
INV_X1M_A9TL40 U76 (.A ( n647 ) , .Y ( n646 ) ) ;
BUF_X1P2M_A9TL40 U75 (.A ( G10 ) , .Y ( n645 ) ) ;
INV_X0P5B_A9TL40 U74 (.A ( G9 ) , .Y ( n644 ) ) ;
INV_X0P7B_A9TL40 U73 (.Y ( n643 ) , .A ( n644 ) ) ;
INV_X0P5B_A9TL40 U72 (.A ( G6 ) , .Y ( n642 ) ) ;
INV_X1B_A9TL40 U71 (.A ( n642 ) , .Y ( n641 ) ) ;
INV_X0P5B_A9TL40 U70 (.A ( G5 ) , .Y ( n640 ) ) ;
INV_X0P8M_A9TL40 U69 (.A ( n640 ) , .Y ( n639 ) ) ;
BUF_X1P2M_A9TL40 U68 (.A ( G4 ) , .Y ( n638 ) ) ;
INV_X0P5B_A9TL40 U67 (.A ( G3 ) , .Y ( n637 ) ) ;
INV_X0P8B_A9TL40 U66 (.A ( n637 ) , .Y ( n636 ) ) ;
INV_X0P5B_A9TL40 U65 (.A ( G2 ) , .Y ( n635 ) ) ;
INV_X0P6M_A9TL40 U64 (.A ( n635 ) , .Y ( n634 ) ) ;
INV_X0P5B_A9TL40 U63 (.A ( G1 ) , .Y ( n633 ) ) ;
INV_X0P6M_A9TL40 U62 (.A ( n633 ) , .Y ( n632 ) ) ;
INV_X0P5B_A9TL40 U61 (.A ( G0 ) , .Y ( n631 ) ) ;
INV_X0P8M_A9TL40 U60 (.A ( n631 ) , .Y ( n630 ) ) ;
INV_X0P5B_A9TL40 U22 (.A ( blif_reset_net ) , .Y ( n629 ) ) ;
INV_X0P5B_A9TL40 U59 (.A ( G13 ) , .Y ( n628 ) ) ;
INV_X1B_A9TL40 U58 (.A ( n628 ) , .Y ( n627 ) ) ;
INV_X0P5B_A9TL40 U57 (.A ( n667 ) , .Y ( n626 ) ) ;
INV_X1M_A9TL40 U56 (.A ( n626 ) , .Y ( n625 ) ) ;
INV_X0P5B_A9TL40 U55 (.A ( n665 ) , .Y ( n624 ) ) ;
INV_X1M_A9TL40 U54 (.A ( n624 ) , .Y ( n623 ) ) ;
INV_X0P5B_A9TL40 U53 (.A ( n663 ) , .Y ( n622 ) ) ;
INV_X1B_A9TL40 U52 (.A ( n622 ) , .Y ( n621 ) ) ;
INV_X0P5B_A9TL40 U51 (.A ( n661 ) , .Y ( n620 ) ) ;
INV_X1M_A9TL40 U50 (.A ( n620 ) , .Y ( n619 ) ) ;
INV_X0P5B_A9TL40 U49 (.A ( G8 ) , .Y ( n618 ) ) ;
INV_X1B_A9TL40 U48 (.A ( n618 ) , .Y ( n617 ) ) ;
INV_X0P5B_A9TL40 U47 (.A ( G7 ) , .Y ( n616 ) ) ;
INV_X0P7B_A9TL40 U46 (.A ( n616 ) , .Y ( n615 ) ) ;
BUF_X1P2M_A9TL40 U45 (.A ( n659 ) , .Y ( n614 ) ) ;
INV_X0P5B_A9TL40 U44 (.A ( n657 ) , .Y ( n613 ) ) ;
INV_X1B_A9TL40 U43 (.A ( n613 ) , .Y ( n612 ) ) ;
INV_X0P5B_A9TL40 U42 (.Y ( n611 ) , .A ( n599 ) ) ;
INV_X1B_A9TL40 U41 (.A ( n611 ) , .Y ( n610 ) ) ;
INV_X0P5B_A9TL40 U40 (.A ( n654 ) , .Y ( n609 ) ) ;
INV_X0P8M_A9TL40 U39 (.A ( n609 ) , .Y ( n608 ) ) ;
INV_X0P5B_A9TL40 U38 (.A ( n652 ) , .Y ( n607 ) ) ;
INV_X0P7B_A9TL40 U37 (.A ( n607 ) , .Y ( n606 ) ) ;
INV_X0P5B_A9TL40 U36 (.A ( n650 ) , .Y ( n605 ) ) ;
INV_X0P8B_A9TL40 U35 (.A ( n605 ) , .Y ( n604 ) ) ;
INV_X0P5B_A9TL40 U24 (.A ( n648 ) , .Y ( n603 ) ) ;
INV_X1M_A9TL40 U23 (.A ( n603 ) , .Y ( n602 ) ) ;
INV_X1B_A9TL40 U4 (.A ( n629 ) , .Y ( n600 ) ) ;
BUF_X1P2M_A9TL40 U3 (.A ( n656 ) , .Y ( n599 ) ) ;
INV_X1B_A9TL40 U34 (.A ( n256 ) , .Y ( n598 ) ) ;
INV_X0P6B_A9TL40 U33 (.A ( n462 ) , .Y ( n597 ) ) ;
INV_X1B_A9TL40 U32 (.A ( n595 ) , .Y ( n596 ) ) ;
BUF_X1P2M_A9TL40 U31 (.A ( n608 ) , .Y ( n595 ) ) ;
INV_X0P8B_A9TL40 U30 (.A ( n593 ) , .Y ( n594 ) ) ;
BUF_X1P2M_A9TL40 U29 (.A ( n606 ) , .Y ( n593 ) ) ;
INV_X0P8B_A9TL40 U28 (.A ( n591 ) , .Y ( n592 ) ) ;
BUFH_X1M_A9TL40 U27 (.A ( n604 ) , .Y ( n591 ) ) ;
INV_X0P5B_A9TL40 U26 (.A ( n589 ) , .Y ( n590 ) ) ;
BUF_X1M_A9TL40 U25 (.A ( n602 ) , .Y ( n589 ) ) ;
INV_X0P8B_A9TL40 U21 (.A ( n584 ) , .Y ( n585 ) ) ;
BUF_X1M_A9TL40 U20 (.A ( n623 ) , .Y ( n584 ) ) ;
INV_X0P8B_A9TL40 U19 (.A ( n582 ) , .Y ( n583 ) ) ;
BUF_X1M_A9TL40 U18 (.A ( n621 ) , .Y ( n582 ) ) ;
INV_X0P8B_A9TL40 U17 (.A ( n580 ) , .Y ( n581 ) ) ;
BUFH_X1M_A9TL40 U16 (.A ( n619 ) , .Y ( n580 ) ) ;
INV_X0P5B_A9TL40 U15 (.A ( n578 ) , .Y ( n579 ) ) ;
BUFH_X1M_A9TL40 U14 (.A ( n617 ) , .Y ( n578 ) ) ;
INV_X0P5B_A9TL40 U13 (.A ( n576 ) , .Y ( n577 ) ) ;
BUF_X1M_A9TL40 U12 (.A ( n615 ) , .Y ( n576 ) ) ;
INV_X1B_A9TL40 U11 (.A ( n574 ) , .Y ( n575 ) ) ;
BUFH_X1M_A9TL40 U10 (.A ( n573 ) , .Y ( n574 ) ) ;
BUF_X1M_A9TL40 U9 (.A ( n614 ) , .Y ( n573 ) ) ;
INV_X0P8B_A9TL40 U8 (.A ( n571 ) , .Y ( n572 ) ) ;
BUFH_X1M_A9TL40 U7 (.A ( n612 ) , .Y ( n571 ) ) ;
INV_X1B_A9TL40 U6 (.A ( n569 ) , .Y ( n570 ) ) ;
BUF_X1M_A9TL40 U5 (.A ( n610 ) , .Y ( n569 ) ) ;
INV_X0P5B_A9TL40 U2 (.A ( n565 ) , .Y ( n566 ) ) ;
BUF_X1M_A9TL40 U1 (.Y ( n565 ) , .A ( n625 ) ) ;
OAI31_X2M_A9TL40 U492 (.B0 ( n434 ) , .A1 ( n490 ) , .Y ( G530 ) , .A0 ( n589 ) 
    , .A2 ( n495 ) ) ;
OAI211_X2M_A9TL40 U568 (.Y ( G551 ) , .A0 ( n505 ) , .A1 ( n504 ) , .B0 ( n503 ) 
    , .C0 ( n502 ) ) ;
AOI22_X1M_A9TL40 U423 (.B0 ( n569 ) , .Y ( n503 ) , .B1 ( n497 ) , .A1 ( n498 ) 
    , .A0 ( n571 ) ) ;
INV_X1M_A9TL40 U302 (.A ( n491 ) , .Y ( n394 ) ) ;
AOI22_X1M_A9TL40 U352 (.B0 ( n470 ) , .Y ( n481 ) , .B1 ( n469 ) , .A1 ( n471 ) 
    , .A0 ( n500 ) ) ;
NOR2_X0P5M_A9TL40 U331 (.B ( n572 ) , .Y ( n492 ) , .A ( n591 ) ) ;
AOI32_X1M_A9TL40 U459 (.A1 ( n580 ) , .A0 ( n441 ) , .A2 ( n312 ) , .Y ( n313 ) 
    , .B0 ( n311 ) , .B1 ( n581 ) ) ;
NAND2_X3B_A9TL40 U533 (.B ( n580 ) , .Y ( n475 ) , .A ( n583 ) ) ;
INV_X0P5B_A9TL40 U332 (.A ( G31 ) , .Y ( n312 ) ) ;
NAND3_X0P5M_A9TL40 U441 (.A ( n565 ) , .Y ( n375 ) , .B ( n359 ) , .C ( n628 ) ) ;
NOR2_X0P5M_A9TL40 U421 (.B ( n583 ) , .Y ( n383 ) , .A ( n579 ) ) ;
NAND2_X0P5M_A9TL40 U471 (.B ( n593 ) , .Y ( n401 ) , .A ( n488 ) ) ;
NAND2_X0P5M_A9TL40 U412 (.B ( n574 ) , .Y ( n297 ) , .A ( n581 ) ) ;
INV_X0P5B_A9TL40 U321 (.A ( n297 ) , .Y ( n449 ) ) ;
INV_X0P5B_A9TL40 U557 (.A ( G34 ) , .Y ( n364 ) ) ;
INV_X0P5B_A9TL40 U320 (.A ( n415 ) , .Y ( n485 ) ) ;
NAND2_X0P5M_A9TL40 U481 (.B ( n593 ) , .Y ( n400 ) , .A ( n569 ) ) ;
NOR3_X0P5M_A9TL40 U411 (.B ( n378 ) , .Y ( n362 ) , .A ( n383 ) , .C ( n577 ) ) ;
NOR3_X0P5M_A9TL40 U417 (.B ( G33 ) , .Y ( n399 ) , .A ( n627 ) , .C ( n596 ) ) ;
OA1B2_X0P5M_A9TL40 U498 (.Y ( n306 ) , .A0N ( n596 ) , .B1 ( n329 ) 
    , .B0 ( n330 ) ) ;
NAND2_X0P5M_A9TL40 U538 (.B ( G30 ) , .Y ( n298 ) , .A ( n576 ) ) ;
NOR2_X0P5M_A9TL40 U489 (.B ( n454 ) , .Y ( n304 ) , .A ( n571 ) ) ;
NOR2_X0P5M_A9TL40 U488 (.B ( n378 ) , .Y ( n301 ) , .A ( n575 ) ) ;
NOR2_X0P5M_A9TL40 U543 (.B ( n256 ) , .Y ( n308 ) , .A ( n414 ) ) ;
NOR3_X0P5M_A9TL40 U496 (.B ( n592 ) , .Y ( n323 ) , .A ( n569 ) , .C ( n359 ) ) ;
NOR3_X0P5M_A9TL40 U497 (.B ( n574 ) , .Y ( n303 ) , .A ( n580 ) , .C ( n453 ) ) ;
NOR3_X0P5M_A9TL40 U303 (.B ( n597 ) , .Y ( n322 ) , .A ( n594 ) , .C ( n345 ) ) ;
INV_X0P5B_A9TL40 U528 (.A ( G41 ) , .Y ( G546 ) ) ;
INV_X0P5B_A9TL40 U299 (.A ( n292 ) , .Y ( n506 ) ) ;
NAND2_X0P5M_A9TL40 U361 (.B ( n482 ) , .Y ( G507 ) , .A ( n394 ) ) ;
NAND2_X0P5M_A9TL40 U544 (.B ( n358 ) , .Y ( G508 ) , .A ( n435 ) ) ;
INV_X0P5B_A9TL40 U545 (.A ( G30 ) , .Y ( n321 ) ) ;
NOR3_X1M_A9TL40 U546 (.B ( n321 ) , .Y ( n310 ) , .A ( n577 ) , .C ( n574 ) ) ;
NOR2_X0P7M_A9TL40 U540 (.B ( n576 ) , .Y ( n332 ) , .A ( n578 ) ) ;
NOR2_X1M_A9TL40 U526 (.B ( n570 ) , .Y ( n462 ) , .A ( n571 ) ) ;
NAND2_X0P5M_A9TL40 U535 (.B ( n576 ) , .Y ( n385 ) , .A ( n582 ) ) ;
NOR2_X1B_A9TL40 U328 (.B ( n575 ) , .Y ( n414 ) , .A ( n570 ) ) ;
NOR2_X0P5M_A9TL40 U530 (.B ( n581 ) , .Y ( n302 ) , .A ( n585 ) ) ;
NOR2_X0P5M_A9TL40 U527 (.B ( n596 ) , .Y ( n487 ) , .A ( n593 ) ) ;
AOI32_X0P7M_A9TL40 U548 (.A1 ( n584 ) , .A0 ( n315 ) , .A2 ( n314 ) 
    , .Y ( n316 ) , .B0 ( n313 ) , .B1 ( n585 ) ) ;
INV_X0P5B_A9TL40 U468 (.A ( n385 ) , .Y ( n423 ) ) ;
INV_X0P5B_A9TL40 U479 (.A ( n475 ) , .Y ( n381 ) ) ;
AOI21_X0P7M_A9TL40 U549 (.B0 ( n316 ) , .Y ( n318 ) , .A1 ( n570 ) 
    , .A0 ( n317 ) ) ;
OAI211_X0P5M_A9TL40 U551 (.Y ( n328 ) , .A0 ( n380 ) , .A1 ( n321 ) 
    , .B0 ( n320 ) , .C0 ( n360 ) ) ;
NOR2_X1B_A9TL40 U461 (.B ( n347 ) , .Y ( n353 ) , .A ( n495 ) ) ;
NAND2_X0P5M_A9TL40 U552 (.B ( G32 ) , .Y ( n345 ) , .A ( n328 ) ) ;
NOR3_X1M_A9TL40 U558 (.B ( n566 ) , .Y ( n428 ) , .A ( n627 ) , .C ( n359 ) ) ;
AOI22_X0P5M_A9TL40 U440 (.B0 ( n491 ) , .Y ( n407 ) , .B1 ( n462 ) 
    , .A1 ( n493 ) , .A0 ( n592 ) ) ;
NAND2_X0P5M_A9TL40 U447 (.B ( n628 ) , .Y ( n369 ) , .A ( n345 ) ) ;
INV_X0P6M_A9TL40 U554 (.A ( n493 ) , .Y ( n482 ) ) ;
AND2_X0P5M_A9TL40 U356 (.B ( n590 ) , .A ( n395 ) , .Y ( n486 ) ) ;
NOR2_X0P5M_A9TL40 U362 (.B ( n418 ) , .Y ( n395 ) , .A ( n499 ) ) ;
NOR2_X1B_A9TL40 U438 (.B ( n482 ) , .Y ( n413 ) , .A ( n592 ) ) ;
NOR2_X1B_A9TL40 U367 (.B ( n369 ) , .Y ( n432 ) , .A ( n371 ) ) ;
NOR2_X0P5M_A9TL40 U297 (.B ( n418 ) , .Y ( n387 ) , .A ( n575 ) ) ;
NOR2_X0P5M_A9TL40 U439 (.B ( n375 ) , .Y ( n451 ) , .A ( n366 ) ) ;
INV_X0P5B_A9TL40 U559 (.A ( n387 ) , .Y ( n426 ) ) ;
NOR2_X0P5M_A9TL40 U360 (.B ( n418 ) , .Y ( n500 ) , .A ( n590 ) ) ;
AOI21_X0P5M_A9TL40 U433 (.B0 ( n405 ) , .Y ( n411 ) , .A1 ( n598 ) 
    , .A0 ( n413 ) ) ;
NAND2_X0P7M_A9TL40 U437 (.B ( n432 ) , .Y ( n438 ) , .A ( n566 ) ) ;
AO21A1AI2_X0P5M_A9TL40 U567 (.B0 ( n490 ) , .Y ( n498 ) , .C0 ( n489 ) 
    , .A1 ( n593 ) , .A0 ( n589 ) ) ;
AOI2XB1_X0P5M_A9TL40 U556 (.A1N ( n432 ) , .A0 ( n439 ) , .Y ( n476 ) 
    , .B0 ( n565 ) ) ;
OA21A1OI2_X0P5M_A9TL40 U560 (.B0 ( n426 ) , .C0 ( n360 ) , .A0 ( n579 ) 
    , .A1 ( n364 ) , .Y ( n422 ) ) ;
NOR2_X0P5M_A9TL40 U565 (.B ( n438 ) , .Y ( n470 ) , .A ( n595 ) ) ;
OAI211_X0P7M_A9TL40 U562 (.Y ( G552 ) , .A0 ( G40 ) , .A1 ( n418 ) 
    , .B0 ( n417 ) , .C0 ( n416 ) ) ;
OA21A1OI2_X0P5M_A9TL40 U566 (.B0 ( n593 ) , .C0 ( n470 ) , .A0 ( n486 ) 
    , .A1 ( n433 ) , .Y ( n434 ) ) ;
NAND2_X0P5B_A9TL40 U476 (.B ( n441 ) , .Y ( n377 ) , .A ( n583 ) ) ;
NOR2_X1M_A9TL40 U477 (.B ( n579 ) , .Y ( n441 ) , .A ( n576 ) ) ;
AND4_X0P5M_A9TL40 U478 (.B ( n570 ) , .C ( n590 ) , .A ( n576 ) , .D ( n583 ) 
    , .Y ( G511 ) ) ;
NAND2_X0P5B_A9TL40 U480 (.B ( n448 ) , .Y ( n406 ) , .A ( n596 ) ) ;
OA21_X0P5M_A9TL40 U482 (.A0 ( n581 ) , .A1 ( n577 ) , .B0 ( n383 ) , .Y ( n420 ) ) ;
NAND2_X0P5B_A9TL40 U483 (.B ( n596 ) , .Y ( n341 ) , .A ( n594 ) ) ;
OAI31_X1M_A9TL40 U485 (.B0 ( n328 ) , .A1 ( n330 ) , .Y ( n368 ) , .A0 ( n331 ) 
    , .A2 ( n329 ) ) ;
NAND3_X0P5M_A9TL40 U486 (.A ( n582 ) , .Y ( n473 ) , .B ( n332 ) , .C ( n302 ) ) ;
NAND3_X0P5M_A9TL40 U490 (.A ( n419 ) , .Y ( n358 ) , .B ( n583 ) , .C ( n575 ) ) ;
OAI22_X0P5M_A9TL40 U491 (.B0 ( n565 ) , .Y ( G539 ) , .A0 ( n376 ) 
    , .A1 ( n375 ) , .B1 ( n374 ) ) ;
OAI22_X0P5M_A9TL40 U493 (.B0 ( n388 ) , .Y ( G547 ) , .A0 ( n389 ) 
    , .A1 ( n426 ) , .B1 ( n581 ) ) ;
NAND3_X0P5M_A9TL40 U494 (.A ( n485 ) , .Y ( n416 ) , .B ( n491 ) , .C ( n597 ) ) ;
NAND3_X0P5M_A9TL40 U495 (.A ( n598 ) , .Y ( n502 ) , .B ( n500 ) , .C ( n499 ) ) ;
OAI22_X0P5M_A9TL40 U499 (.B0 ( n390 ) , .Y ( n307 ) , .A0 ( n592 ) 
    , .A1 ( n415 ) , .B1 ( n429 ) ) ;
OAI31_X0P5M_A9TL40 U500 (.B0 ( n295 ) , .A1 ( n574 ) , .Y ( n296 ) 
    , .A0 ( n381 ) , .A2 ( n577 ) ) ;
AO21A1AI2_X0P5M_A9TL40 U501 (.B0 ( n300 ) , .Y ( G513 ) , .C0 ( n578 ) 
    , .A1 ( n583 ) , .A0 ( n301 ) ) ;
AOI21_X0P5M_A9TL40 U502 (.B0 ( n294 ) , .Y ( G502 ) , .A1 ( n597 ) 
    , .A0 ( n487 ) ) ;
NAND3_X0P5M_A9TL40 U503 (.A ( n593 ) , .Y ( n293 ) , .B ( n492 ) , .C ( n570 ) ) ;
OA21_X0P5M_A9TL40 U523 (.A0 ( n580 ) , .A1 ( n585 ) , .B0 ( n583 ) , .Y ( n287 ) ) ;
NAND3_X0P5M_A9TL40 U524 (.A ( n591 ) , .Y ( n490 ) , .B ( n428 ) , .C ( n596 ) ) ;
AO21A1AI2_X0P5M_A9TL40 U525 (.B0 ( n590 ) , .Y ( n291 ) , .C0 ( n591 ) 
    , .A1 ( n570 ) , .A0 ( n595 ) ) ;
OAI21_X0P5M_A9TL40 U529 (.A0 ( n574 ) , .A1 ( n581 ) , .Y ( G510 ) 
    , .B0 ( n297 ) ) ;
OAI22_X0P5M_A9TL40 U531 (.B0 ( n302 ) , .Y ( G504 ) , .A0 ( n576 ) 
    , .A1 ( n585 ) , .B1 ( n583 ) ) ;
AOI22_X0P5M_A9TL40 U532 (.B0 ( n256 ) , .Y ( G512 ) , .B1 ( n594 ) 
    , .A1 ( n598 ) , .A0 ( n593 ) ) ;
AOI21_X0P5M_A9TL40 U534 (.B0 ( n419 ) , .Y ( n295 ) , .A1 ( n449 ) 
    , .A0 ( n383 ) ) ;
AOI22_X0P5M_A9TL40 U536 (.B0 ( n301 ) , .Y ( G515 ) , .B1 ( n385 ) 
    , .A1 ( n296 ) , .A0 ( n584 ) ) ;
OAI211_X0P5M_A9TL40 U537 (.Y ( n299 ) , .A0 ( n575 ) , .A1 ( n585 ) 
    , .B0 ( n576 ) , .C0 ( n297 ) ) ;
AOI22_X0P5M_A9TL40 U539 (.B0 ( n575 ) , .Y ( n300 ) , .B1 ( n298 ) 
    , .A1 ( n299 ) , .A0 ( n312 ) ) ;
NAND2XB_X0P5M_A9TL40 U541 (.A ( n453 ) , .Y ( G509 ) , .BN ( n304 ) ) ;
NAND2_X1M_A9TL40 U542 (.B ( n593 ) , .Y ( n495 ) , .A ( n571 ) ) ;
AOI211_X1M_A9TL40 U547 (.B0 ( n582 ) , .Y ( n311 ) , .C0 ( n310 ) , .A1 ( G31 ) 
    , .A0 ( n578 ) ) ;
OAI211_X1M_A9TL40 U550 (.Y ( n359 ) , .A0 ( n338 ) , .A1 ( n319 ) , .B0 ( G46 ) 
    , .C0 ( n318 ) ) ;
NOR3_X1A_A9TL40 U553 (.B ( n627 ) , .Y ( n491 ) , .A ( n565 ) , .C ( n345 ) ) ;
NAND2_X0P5B_A9TL40 U555 (.B ( n627 ) , .Y ( n439 ) , .A ( n367 ) ) ;
OAI22_X0P5M_A9TL40 U561 (.B0 ( G42 ) , .Y ( G548 ) , .A0 ( n365 ) , .A1 ( n364 ) 
    , .B1 ( n418 ) ) ;
OAI21_X0P5M_A9TL40 U563 (.A0 ( n578 ) , .A1 ( n585 ) , .Y ( n421 ) 
    , .B0 ( n580 ) ) ;
NAND2_X0P5B_A9TL40 U564 (.B ( n598 ) , .Y ( n430 ) , .A ( n570 ) ) ;
NAND2_X0P5B_A9TL40 U383 (.B ( n574 ) , .Y ( n435 ) , .A ( n336 ) ) ;
NAND2XB_X0P5M_A9TL40 U384 (.A ( n353 ) , .Y ( n445 ) , .BN ( n454 ) ) ;
AOI211_X0P5M_A9TL40 U385 (.B0 ( n484 ) , .Y ( n505 ) , .C0 ( n483 ) 
    , .A1 ( n572 ) , .A0 ( n485 ) ) ;
AO21A1AI2_X0P5M_A9TL40 U386 (.B0 ( n484 ) , .Y ( n288 ) , .C0 ( n589 ) 
    , .A1 ( n597 ) , .A0 ( n341 ) ) ;
AOI21_X0P5M_A9TL40 U387 (.B0 ( n325 ) , .Y ( n327 ) , .A1 ( n390 ) 
    , .A0 ( n598 ) ) ;
AOI22_X0P5M_A9TL40 U388 (.B0 ( G36 ) , .Y ( n342 ) , .B1 ( n575 ) , .A1 ( n336 ) 
    , .A0 ( n467 ) ) ;
NAND2_X0P5B_A9TL40 U389 (.B ( n346 ) , .Y ( n472 ) , .A ( n572 ) ) ;
NOR3_X0P7M_A9TL40 U390 (.B ( n585 ) , .Y ( n467 ) , .A ( n572 ) , .C ( n390 ) ) ;
AOI21_X0P5M_A9TL40 U391 (.B0 ( n362 ) , .Y ( n365 ) , .A1 ( n363 ) 
    , .A0 ( n584 ) ) ;
OAI22BB_X0P5M_A9TL40 U392 (.A0 ( n594 ) , .A1 ( n597 ) , .Y ( n393 ) 
    , .B1N ( n487 ) , .B0N ( n571 ) ) ;
AOI21_X0P5M_A9TL40 U393 (.B0 ( n379 ) , .Y ( n389 ) , .A1 ( n380 ) 
    , .A0 ( n381 ) ) ;
OAI31_X0P5M_A9TL40 U394 (.B0 ( n333 ) , .A1 ( n406 ) , .Y ( n335 ) 
    , .A0 ( n571 ) , .A2 ( n334 ) ) ;
NOR3_X0P7M_A9TL40 U395 (.B ( n499 ) , .Y ( n330 ) , .A ( n574 ) , .C ( n594 ) ) ;
OAI22_X0P5M_A9TL40 U396 (.B0 ( n465 ) , .Y ( n348 ) , .A0 ( n591 ) 
    , .A1 ( n347 ) , .B1 ( n410 ) ) ;
OAI22_X0P5M_A9TL40 U397 (.B0 ( n571 ) , .Y ( n402 ) , .A0 ( n488 ) 
    , .A1 ( n495 ) , .B1 ( n401 ) ) ;
OAI211_X0P5M_A9TL40 U398 (.Y ( n384 ) , .A0 ( n576 ) , .A1 ( n383 ) 
    , .B0 ( G34 ) , .C0 ( n382 ) ) ;
NAND3_X0P7M_A9TL40 U399 (.A ( n578 ) , .Y ( n454 ) , .B ( n423 ) , .C ( n302 ) ) ;
OAI21_X0P5M_A9TL40 U400 (.A0 ( n579 ) , .A1 ( n378 ) , .Y ( n320 ) 
    , .B0 ( n423 ) ) ;
NAND2_X0P5B_A9TL40 U401 (.B ( n414 ) , .Y ( n347 ) , .A ( n595 ) ) ;
OAI22_X0P5M_A9TL40 U402 (.B0 ( n580 ) , .Y ( n363 ) , .A0 ( n381 ) 
    , .A1 ( n380 ) , .B1 ( n385 ) ) ;
AOI21_X0P5M_A9TL40 U403 (.B0 ( n462 ) , .Y ( n324 ) , .A1 ( n574 ) 
    , .A0 ( n593 ) ) ;
NAND3B_X0P5M_A9TL40 U404 (.C ( n583 ) , .AN ( n338 ) , .B ( n572 ) , .Y ( n453 ) ) ;
AOI22_X0P5M_A9TL40 U405 (.B0 ( n575 ) , .Y ( n315 ) , .B1 ( n321 ) 
    , .A1 ( n581 ) , .A0 ( n332 ) ) ;
AOI211_X0P5M_A9TL40 U406 (.B0 ( n420 ) , .Y ( n427 ) , .C0 ( n419 ) 
    , .A1 ( n421 ) , .A0 ( n582 ) ) ;
AOI21_X0P5M_A9TL40 U407 (.B0 ( n492 ) , .Y ( n431 ) , .A1 ( n256 ) 
    , .A0 ( n569 ) ) ;
NAND2_X0P5B_A9TL40 U408 (.B ( n575 ) , .Y ( n466 ) , .A ( n570 ) ) ;
OR2_X0P5M_A9TL40 U409 (.Y ( n429 ) , .B ( n571 ) , .A ( n465 ) ) ;
NAND2_X0P5B_A9TL40 U410 (.B ( n332 ) , .Y ( n338 ) , .A ( n585 ) ) ;
NAND4_X0P7M_A9TL40 U413 (.C ( n572 ) , .B ( n337 ) , .D ( n570 ) , .Y ( n436 ) 
    , .A ( n595 ) ) ;
NAND2_X0P5B_A9TL40 U414 (.B ( n595 ) , .Y ( n465 ) , .A ( n591 ) ) ;
NOR3_X0P7M_A9TL40 U415 (.B ( n580 ) , .Y ( n419 ) , .A ( n578 ) , .C ( n577 ) ) ;
NAND2_X0P5B_A9TL40 U416 (.B ( n576 ) , .Y ( n309 ) , .A ( n581 ) ) ;
NAND2_X0P5B_A9TL40 U418 (.B ( n580 ) , .Y ( n319 ) , .A ( n582 ) ) ;
NOR2_X0P7M_A9TL40 U419 (.B ( n575 ) , .Y ( n448 ) , .A ( n569 ) ) ;
AOI22_X0P5M_A9TL40 U420 (.B0 ( n571 ) , .Y ( n317 ) , .B1 ( n596 ) 
    , .A1 ( n589 ) , .A0 ( n595 ) ) ;
OAI211_X0P7M_A9TL40 U422 (.Y ( G542 ) , .A0 ( n427 ) , .A1 ( n426 ) 
    , .B0 ( n425 ) , .C0 ( n424 ) ) ;
AOI31_X0P7M_A9TL40 U424 (.A1 ( n413 ) , .A0 ( n414 ) , .Y ( n417 ) 
    , .A2 ( n495 ) , .B0 ( n412 ) ) ;
OAI211_X0P7M_A9TL40 U425 (.Y ( G550 ) , .A0 ( G29 ) , .A1 ( n496 ) 
    , .B0 ( n404 ) , .C0 ( n403 ) ) ;
OAI211_X0P5M_A9TL40 U426 (.Y ( G549 ) , .A0 ( n398 ) , .A1 ( n504 ) 
    , .B0 ( n397 ) , .C0 ( n396 ) ) ;
OAI211_X0P5M_A9TL40 U427 (.Y ( G532 ) , .A0 ( G43 ) , .A1 ( n482 ) 
    , .B0 ( n481 ) , .C0 ( n480 ) ) ;
AOI31_X0P7M_A9TL40 U428 (.A1 ( n430 ) , .A0 ( n431 ) , .Y ( n433 ) 
    , .A2 ( n429 ) , .B0 ( n496 ) ) ;
OAI31_X0P7M_A9TL40 U429 (.B0 ( n494 ) , .A1 ( n496 ) , .Y ( n497 ) 
    , .A0 ( n595 ) , .A2 ( n495 ) ) ;
OAI22_X0P7M_A9TL40 U430 (.B0 ( n409 ) , .Y ( n412 ) , .A0 ( n411 ) 
    , .A1 ( n410 ) , .B1 ( n594 ) ) ;
AOI211_X0P7M_A9TL40 U431 (.B0 ( n399 ) , .Y ( n397 ) , .C0 ( n486 ) 
    , .A1 ( n570 ) , .A0 ( n405 ) ) ;
OAI31_X0P5M_A9TL40 U432 (.B0 ( n476 ) , .A1 ( n478 ) , .Y ( n480 ) 
    , .A0 ( n479 ) , .A2 ( n477 ) ) ;
NOR2XB_X0P7M_A9TL40 U434 (.Y ( n450 ) , .A ( n437 ) , .BN ( G38 ) ) ;
OAI31_X0P7M_A9TL40 U435 (.B0 ( n384 ) , .A1 ( n418 ) , .Y ( n386 ) 
    , .A0 ( n574 ) , .A2 ( n385 ) ) ;
OAI22_X0P7M_A9TL40 U436 (.B0 ( n482 ) , .Y ( n408 ) , .A0 ( n575 ) 
    , .A1 ( n407 ) , .B1 ( n406 ) ) ;
INV_X0P6B_A9TL40 U442 (.A ( n369 ) , .Y ( n370 ) ) ;
NOR2XB_X0P5M_A9TL40 U443 (.Y ( n372 ) , .A ( n628 ) , .BN ( n368 ) ) ;
NOR3_X2M_A9TL40 U444 (.A ( n565 ) , .Y ( n493 ) , .B ( n628 ) , .C ( n368 ) ) ;
OAI211_X0P7M_A9TL40 U445 (.Y ( n343 ) , .A0 ( n342 ) , .A1 ( n341 ) 
    , .B0 ( n340 ) , .C0 ( n445 ) ) ;
OAI31_X0P5M_A9TL40 U446 (.B0 ( n289 ) , .A1 ( n574 ) , .Y ( n290 ) 
    , .A0 ( n582 ) , .A2 ( G30 ) ) ;
AO21A1AI2_X0P7M_A9TL40 U448 (.B0 ( n452 ) , .Y ( n366 ) , .C0 ( n591 ) 
    , .A1 ( n335 ) , .A0 ( n337 ) ) ;
OAI31_X0P5M_A9TL40 U449 (.B0 ( n350 ) , .A1 ( n378 ) , .Y ( n356 ) 
    , .A0 ( n351 ) , .A2 ( n377 ) ) ;
OA21A1OI2_X0P7M_A9TL40 U450 (.B0 ( n446 ) , .C0 ( n472 ) , .A0 ( n380 ) 
    , .A1 ( n475 ) , .Y ( n344 ) ) ;
OAI21_X0P5M_A9TL40 U451 (.A0 ( n446 ) , .A1 ( n472 ) , .Y ( n447 ) 
    , .B0 ( n445 ) ) ;
AOI31_X0P7M_A9TL40 U452 (.A1 ( n415 ) , .A0 ( n327 ) , .Y ( n331 ) 
    , .A2 ( n391 ) , .B0 ( n592 ) ) ;
AOI211_X0P7M_A9TL40 U453 (.B0 ( n592 ) , .Y ( n355 ) , .C0 ( n474 ) 
    , .A1 ( n354 ) , .A0 ( n454 ) ) ;
NAND2_X0P5B_A9TL40 U454 (.B ( n346 ) , .Y ( n351 ) , .A ( n592 ) ) ;
OAI22_X0P5M_A9TL40 U455 (.B0 ( n466 ) , .Y ( n456 ) , .A0 ( n597 ) 
    , .A1 ( n454 ) , .B1 ( n453 ) ) ;
OAI211_X0P5M_A9TL40 U456 (.Y ( n392 ) , .A0 ( n569 ) , .A1 ( n256 ) 
    , .B0 ( n406 ) , .C0 ( n391 ) ) ;
AO21B_X0P5M_A9TL40 U457 (.A0 ( n468 ) , .A1 ( n467 ) , .Y ( n469 ) 
    , .B0N ( n466 ) ) ;
AO21A1AI2_X0P5M_A9TL40 U458 (.B0 ( n349 ) , .Y ( n350 ) , .C0 ( n348 ) 
    , .A1 ( n468 ) , .A0 ( n584 ) ) ;
OAI211_X0P5M_A9TL40 U460 (.Y ( n471 ) , .A0 ( n569 ) , .A1 ( n465 ) 
    , .B0 ( n464 ) , .C0 ( n463 ) ) ;
NAND2_X0P5B_A9TL40 U462 (.B ( n326 ) , .Y ( n391 ) , .A ( n571 ) ) ;
NAND2_X0P5B_A9TL40 U463 (.B ( n423 ) , .Y ( n382 ) , .A ( n578 ) ) ;
OAI211_X0P5M_A9TL40 U464 (.Y ( n424 ) , .A0 ( n579 ) , .A1 ( n581 ) 
    , .B0 ( n423 ) , .C0 ( G34 ) ) ;
INV_X0P6B_A9TL40 U465 (.A ( n473 ) , .Y ( n349 ) ) ;
OAI22_X0P5M_A9TL40 U466 (.B0 ( n585 ) , .Y ( n379 ) , .A0 ( n578 ) 
    , .A1 ( n378 ) , .B1 ( n377 ) ) ;
AO21A1AI2_X0P5M_A9TL40 U467 (.B0 ( n462 ) , .Y ( n464 ) , .C0 ( n596 ) 
    , .A1 ( n594 ) , .A0 ( n591 ) ) ;
OAI31_X0P5M_A9TL40 U469 (.B0 ( n293 ) , .A1 ( n596 ) , .Y ( n294 ) 
    , .A0 ( n591 ) , .A2 ( n400 ) ) ;
NAND2_X0P7B_A9TL40 U470 (.B ( n576 ) , .Y ( n360 ) , .A ( n381 ) ) ;
NAND4XXXB_X1M_A9TL40 U472 (.DN ( n310 ) , .A ( n578 ) , .Y ( n314 ) 
    , .B ( n312 ) , .C ( n475 ) ) ;
AOI211_X0P7M_A9TL40 U473 (.B0 ( n591 ) , .Y ( n329 ) , .C0 ( n594 ) 
    , .A1 ( n410 ) , .A0 ( n572 ) ) ;
NAND4_X0P5A_A9TL40 U474 (.C ( n590 ) , .B ( n332 ) , .D ( n581 ) , .Y ( n334 ) 
    , .A ( n582 ) ) ;
OAI221_X0P5M_A9TL40 U475 (.B1 ( n465 ) , .B0 ( n594 ) , .A1 ( n598 ) 
    , .A0 ( n593 ) , .Y ( n463 ) , .C0 ( n569 ) ) ;
INV_X0P6B_A9TL40 U290 (.A ( n422 ) , .Y ( n425 ) ) ;
AOI211_X0P5M_A9TL40 U291 (.B0 ( n422 ) , .Y ( G514 ) , .C0 ( n361 ) 
    , .A1 ( n420 ) , .A0 ( G34 ) ) ;
INV_X0P6B_A9TL40 U292 (.A ( n476 ) , .Y ( n460 ) ) ;
AOI21_X0P5M_A9TL40 U293 (.B0 ( n408 ) , .Y ( n409 ) , .A1 ( n491 ) 
    , .A0 ( n483 ) ) ;
INV_X0P7B_A9TL40 U294 (.A ( n413 ) , .Y ( n504 ) ) ;
INV_X0P6B_A9TL40 U295 (.A ( n470 ) , .Y ( n444 ) ) ;
INV_X0P7B_A9TL40 U296 (.A ( n500 ) , .Y ( n496 ) ) ;
OAI22_X0P5M_A9TL40 U298 (.B0 ( n438 ) , .Y ( n440 ) , .A0 ( n565 ) 
    , .A1 ( n439 ) , .B1 ( n472 ) ) ;
INV_X0P6B_A9TL40 U300 (.A ( n366 ) , .Y ( n376 ) ) ;
OAI31_X1M_A9TL40 U301 (.B0 ( n357 ) , .A1 ( n436 ) , .Y ( n367 ) , .A0 ( n591 ) 
    , .A2 ( n358 ) ) ;
NOR2_X0P7M_A9TL40 U304 (.B ( n435 ) , .Y ( n479 ) , .A ( n436 ) ) ;
INV_X0P6B_A9TL40 U305 (.A ( n353 ) , .Y ( n474 ) ) ;
INV_X0P7B_A9TL40 U306 (.A ( n446 ) , .Y ( n336 ) ) ;
NOR2_X0P5A_A9TL40 U307 (.B ( n597 ) , .Y ( n484 ) , .A ( n487 ) ) ;
INV_X0P6B_A9TL40 U308 (.A ( n352 ) , .Y ( n354 ) ) ;
NOR2_X0P7M_A9TL40 U309 (.B ( n390 ) , .Y ( n483 ) , .A ( n595 ) ) ;
NOR3_X0P5A_A9TL40 U310 (.B ( n390 ) , .Y ( n457 ) , .A ( n572 ) , .C ( n473 ) ) ;
OAI22_X0P5M_A9TL40 U311 (.B0 ( n595 ) , .Y ( n325 ) , .A0 ( n598 ) 
    , .A1 ( n390 ) , .B1 ( n324 ) ) ;
INV_X0P7B_A9TL40 U312 (.A ( n347 ) , .Y ( n346 ) ) ;
AOI2XB1_X0P5M_A9TL40 U313 (.A1N ( n319 ) , .A0 ( n332 ) , .Y ( n446 ) 
    , .B0 ( n468 ) ) ;
NOR2_X0P7M_A9TL40 U314 (.B ( n338 ) , .Y ( n352 ) , .A ( n475 ) ) ;
INV_X0P7B_A9TL40 U315 (.A ( n436 ) , .Y ( n339 ) ) ;
INV_X0P7B_A9TL40 U316 (.A ( n488 ) , .Y ( n499 ) ) ;
NAND4_X0P5A_A9TL40 U317 (.C ( G37 ) , .B ( n598 ) , .D ( G511 ) , .Y ( n333 ) 
    , .A ( n578 ) ) ;
INV_X0P7B_A9TL40 U319 (.A ( n414 ) , .Y ( n390 ) ) ;
INV_X0P7B_A9TL40 U322 (.A ( n466 ) , .Y ( n326 ) ) ;
NOR2_X1B_A9TL40 U323 (.B ( n592 ) , .Y ( n488 ) , .A ( n570 ) ) ;
NAND2_X0P5B_A9TL40 U324 (.B ( n487 ) , .Y ( n415 ) , .A ( n574 ) ) ;
INV_X0P7B_A9TL40 U325 (.A ( n448 ) , .Y ( n410 ) ) ;
NOR3_X1M_A9TL40 U326 (.B ( n579 ) , .Y ( n468 ) , .A ( n582 ) , .C ( n309 ) ) ;
INV_X0P7B_A9TL40 U327 (.A ( n441 ) , .Y ( n380 ) ) ;
INV_X0P7B_A9TL40 U330 (.A ( n302 ) , .Y ( n378 ) ) ;
NOR2_X0P5A_A9TL40 U337 (.B ( n594 ) , .Y ( n337 ) , .A ( n585 ) ) ;
OR2_X0P7M_A9TL40 U343 (.Y ( n256 ) , .B ( n596 ) , .A ( n572 ) ) ;
OAI211_X0P5M_A9TL40 U344 (.Y ( G535 ) , .A0 ( G44 ) , .A1 ( n444 ) 
    , .B0 ( n443 ) , .C0 ( n442 ) ) ;
OAI211_X0P5M_A9TL40 U345 (.Y ( G537 ) , .A0 ( n461 ) , .A1 ( n460 ) 
    , .B0 ( n459 ) , .C0 ( n458 ) ) ;
AOI22_X0P5M_A9TL40 U346 (.B0 ( n493 ) , .Y ( n403 ) , .B1 ( n402 ) 
    , .A1 ( n486 ) , .A0 ( n595 ) ) ;
AOI22_X0P5M_A9TL40 U347 (.B0 ( G37 ) , .Y ( n443 ) , .B1 ( n450 ) , .A1 ( n479 ) 
    , .A0 ( n476 ) ) ;
AOI31_X0P5M_A9TL40 U348 (.A1 ( n487 ) , .A0 ( n488 ) , .A2 ( n493 ) 
    , .Y ( n489 ) , .B0 ( n486 ) ) ;
AOI22_X0P5M_A9TL40 U349 (.B0 ( n450 ) , .Y ( n459 ) , .B1 ( n449 ) 
    , .A1 ( n451 ) , .A0 ( n452 ) ) ;
NAND2XB_X0P5M_A9TL40 U350 (.A ( n460 ) , .Y ( G518 ) , .BN ( n451 ) ) ;
OAI21_X0P5M_A9TL40 U351 (.A0 ( n441 ) , .A1 ( n468 ) , .Y ( n442 ) 
    , .B0 ( n440 ) ) ;
OAI21_X0P5M_A9TL40 U353 (.A0 ( n457 ) , .A1 ( n456 ) , .Y ( n458 ) 
    , .B0 ( n470 ) ) ;
AOI31_X0P5M_A9TL40 U354 (.A1 ( n441 ) , .A0 ( n582 ) , .A2 ( n387 ) 
    , .Y ( n388 ) , .B0 ( n386 ) ) ;
OAI21_X0P5M_A9TL40 U355 (.A0 ( n395 ) , .A1 ( n405 ) , .Y ( n396 ) 
    , .B0 ( n596 ) ) ;
NAND2_X0P5B_A9TL40 U357 (.B ( n451 ) , .Y ( n437 ) , .A ( n598 ) ) ;
AOI211_X0P5M_A9TL40 U358 (.B0 ( n418 ) , .Y ( n361 ) , .C0 ( n385 ) 
    , .A1 ( n574 ) , .A0 ( n580 ) ) ;
AOI22_X0P5M_A9TL40 U359 (.B0 ( n371 ) , .Y ( n374 ) , .B1 ( n370 ) 
    , .A1 ( n372 ) , .A0 ( n373 ) ) ;
INV_X0P6B_A9TL40 U363 (.A ( n367 ) , .Y ( n373 ) ) ;
AOI32_X0P5M_A9TL40 U364 (.A1 ( n565 ) , .A0 ( n589 ) , .A2 ( n323 ) 
    , .Y ( G506 ) , .B0 ( n322 ) , .B1 ( n566 ) ) ;
AOI22_X0P5M_A9TL40 U365 (.B0 ( n491 ) , .Y ( n494 ) , .B1 ( G39 ) , .A1 ( n492 ) 
    , .A0 ( n493 ) ) ;
AOI31_X0P5M_A9TL40 U366 (.A1 ( n431 ) , .A0 ( n593 ) , .A2 ( n291 ) 
    , .Y ( n292 ) , .B0 ( n290 ) ) ;
NOR2_X1B_A9TL40 U368 (.B ( n394 ) , .Y ( n405 ) , .A ( n495 ) ) ;
AOI31_X1M_A9TL40 U369 (.A1 ( n344 ) , .A0 ( n584 ) , .A2 ( n594 ) , .Y ( n371 ) 
    , .B0 ( n343 ) ) ;
AOI21_X0P5M_A9TL40 U370 (.B0 ( n447 ) , .Y ( n461 ) , .A1 ( n468 ) 
    , .A0 ( n448 ) ) ;
AOI31_X0P5M_A9TL40 U371 (.A1 ( n598 ) , .A0 ( n491 ) , .A2 ( n400 ) 
    , .Y ( n404 ) , .B0 ( n399 ) ) ;
AOI31_X0P5M_A9TL40 U372 (.A1 ( n572 ) , .A0 ( n593 ) , .A2 ( n356 ) 
    , .Y ( n357 ) , .B0 ( n355 ) ) ;
AOI22_X0P5M_A9TL40 U373 (.B0 ( n575 ) , .Y ( n289 ) , .B1 ( n577 ) 
    , .A1 ( n288 ) , .A0 ( n592 ) ) ;
AOI211_X0P5M_A9TL40 U374 (.B0 ( n307 ) , .Y ( G516 ) , .C0 ( n306 ) 
    , .A1 ( n308 ) , .A0 ( n591 ) ) ;
AOI211_X0P5M_A9TL40 U375 (.B0 ( n393 ) , .Y ( n398 ) , .C0 ( n392 ) 
    , .A1 ( n483 ) , .A0 ( n571 ) ) ;
NOR2_X0P5A_A9TL40 U376 (.B ( n472 ) , .Y ( n478 ) , .A ( n473 ) ) ;
OAI21_X0P5M_A9TL40 U377 (.A0 ( n346 ) , .A1 ( n495 ) , .Y ( G505 ) 
    , .B0 ( n305 ) ) ;
NOR2_X0P7M_A9TL40 U378 (.B ( n445 ) , .Y ( n452 ) , .A ( n590 ) ) ;
NOR2_X0P5A_A9TL40 U379 (.B ( n474 ) , .Y ( n477 ) , .A ( n475 ) ) ;
AOI211_X0P5M_A9TL40 U380 (.B0 ( n457 ) , .Y ( G517 ) , .C0 ( n303 ) 
    , .A1 ( n304 ) , .A0 ( n326 ) ) ;
AOI22_X0P5M_A9TL40 U381 (.B0 ( n352 ) , .Y ( n340 ) , .B1 ( n353 ) , .A1 ( G35 ) 
    , .A0 ( n339 ) ) ;
AOI21_X0P5M_A9TL40 U382 (.B0 ( n393 ) , .Y ( n305 ) , .A1 ( n448 ) 
    , .A0 ( n487 ) ) ;
DFFRPQ_X0P5M_A9TL40 G29_reg (.Q ( G29 ) , .CK ( blif_clk_net ) , .D ( G502 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G31_reg (.Q ( G31 ) , .CK ( blif_clk_net ) , .D ( G504 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G32_reg (.Q ( G32 ) , .CK ( blif_clk_net ) , .D ( G505 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G34_reg (.Q ( G34 ) , .CK ( blif_clk_net ) , .D ( G507 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G35_reg (.Q ( G35 ) , .CK ( blif_clk_net ) , .D ( G508 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G36_reg (.Q ( G36 ) , .CK ( blif_clk_net ) , .D ( G509 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G37_reg (.Q ( G37 ) , .CK ( blif_clk_net ) , .D ( G510 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G38_reg (.Q ( G38 ) , .CK ( blif_clk_net ) , .D ( G511 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G39_reg (.Q ( G39 ) , .CK ( blif_clk_net ) , .D ( G512 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G40_reg (.Q ( G40 ) , .CK ( blif_clk_net ) , .D ( G513 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G42_reg (.Q ( G42 ) , .CK ( blif_clk_net ) , .D ( G515 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G43_reg (.Q ( G43 ) , .CK ( blif_clk_net ) , .D ( G516 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G44_reg (.Q ( G44 ) , .CK ( blif_clk_net ) , .D ( G517 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G33_reg (.Q ( G33 ) , .CK ( blif_clk_net ) , .D ( G506 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G41_reg (.Q ( G41 ) , .CK ( blif_clk_net ) , .D ( G514 ) 
    , .R ( n600 ) ) ;
DFFRPQ_X0P5M_A9TL40 G45_reg (.Q ( G45 ) , .CK ( blif_clk_net ) , .D ( G518 ) 
    , .R ( n600 ) ) ;
DFFSQN_X0P5M_A9TL40 G46_reg (.QN ( G46 ) , .D ( n506 ) , .CK ( blif_clk_net ) 
    , .SN ( n629 ) ) ;
DFFSQN_X0P5M_A9TL40 G30_reg (.QN ( G30 ) , .D ( n287 ) , .CK ( blif_clk_net ) 
    , .SN ( n629 ) ) ;
INV_X1B_A9TL40 U289 (.A ( n428 ) , .Y ( n418 ) ) ;
endmodule

