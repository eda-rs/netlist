module s1238_bench
(blif_reset_net  , blif_clk_net  , G548  , G3  , G11  , G2  , G0  , G535  , G6  , G12  , G9  , G539  , G542  , G45  , G530  , G13  , G5  , G551  , G537  , G7  , G1  , G4  , G546  , G547  , G552  , G532  , G549  , G550  , G8  , G10 );
input G3 ;
input G2 ;
input G1 ;
input G0 ;
input blif_reset_net ;
input blif_clk_net ;
input G11 ;
input G10 ;
input G9 ;
input G8 ;
input G7 ;
input G6 ;
input G5 ;
input G4 ;
output G546 ;
output G542 ;
output G552 ;
output G551 ;
output G550 ;
output G549 ;
input G13 ;
input G12 ;
output G539 ;
output G45 ;
output G537 ;
output G535 ;
output G532 ;
output G530 ;
output G548 ;
output G547 ;
INV_X1M_A9TL40 U76  (.Y ( n646 ));
INV_X0P8M_A9TL40 U97  (.A ( n668 ) , .Y ( n667 ));
INV_X0P5B_A9TL40 U57  (.A ( n667 ) , .Y ( n626 ));
INV_X1M_A9TL40 U95  (.A ( n666 ) , .Y ( n665 ));
INV_X0P5B_A9TL40 U55  (.A ( n665 ) , .Y ( n624 ));
BUF_X1P2M_A9TL40 U75  (.Y ( n645 ) , .A ( G10 ));
INV_X0P6M_A9TL40 U93  (.A ( n664 ) , .Y ( n663 ));
INV_X0P5B_A9TL40 U53  (.A ( n663 ) , .Y ( n622 ));
INV_X0P7B_A9TL40 U73  (.Y ( n643 ));
INV_X0P6M_A9TL40 U91  (.A ( n662 ) , .Y ( n661 ));
INV_X0P5B_A9TL40 U51  (.A ( n661 ) , .Y ( n620 ));
INV_X1B_A9TL40 U71  (.Y ( n641 ));
INV_X1B_A9TL40 U89  (.A ( n660 ) , .Y ( n659 ));
BUF_X1P2M_A9TL40 U45  (.A ( n659 ) , .Y ( n614 ));
INV_X0P8M_A9TL40 U69  (.Y ( n639 ));
INV_X0P8M_A9TL40 U87  (.A ( n658 ) , .Y ( n657 ));
INV_X0P5B_A9TL40 U44  (.A ( n657 ) , .Y ( n613 ));
BUF_X1P2M_A9TL40 U68  (.Y ( n638 ) , .A ( G4 ));
BUF_X1P2M_A9TL40 U3  (.A ( n656 ));
INV_X0P8B_A9TL40 U66  (.Y ( n636 ));
INV_X0P7B_A9TL40 U84  (.A ( n655 ) , .Y ( n654 ));
INV_X0P5B_A9TL40 U40  (.A ( n654 ) , .Y ( n609 ));
INV_X0P6M_A9TL40 U64  (.Y ( n634 ));
INV_X0P7B_A9TL40 U82  (.A ( n653 ) , .Y ( n652 ));
INV_X0P5B_A9TL40 U38  (.A ( n652 ) , .Y ( n607 ));
INV_X0P6M_A9TL40 U62  (.Y ( n632 ));
INV_X0P7B_A9TL40 U80  (.A ( n651 ) , .Y ( n650 ));
INV_X0P5B_A9TL40 U36  (.A ( n650 ) , .Y ( n605 ));
INV_X0P8M_A9TL40 U60  (.Y ( n630 ));
INV_X0P8M_A9TL40 U78  (.A ( n649 ) , .Y ( n648 ));
INV_X0P5B_A9TL40 U24  (.A ( n648 ) , .Y ( n603 ));
INV_X1M_A9TL40 U76  (.A ( n647 ));
INV_X0P7B_A9TL40 U73  (.A ( n644 ));
INV_X1B_A9TL40 U71  (.A ( n642 ));
INV_X0P8M_A9TL40 U69  (.A ( n640 ));
INV_X0P8B_A9TL40 U66  (.A ( n637 ));
INV_X0P6M_A9TL40 U64  (.A ( n635 ));
INV_X0P6M_A9TL40 U62  (.A ( n633 ));
INV_X0P8M_A9TL40 U60  (.A ( n631 ));
INV_X1B_A9TL40 U4  (.A ( n629 ) , .Y ( n600 ));
DFFSQN_X0P5M_A9TL40 G46_reg  (.SN ( n629 ));
DFFSQN_X0P5M_A9TL40 G30_reg  (.SN ( n629 ));
INV_X1B_A9TL40 U58  (.A ( n628 ) , .Y ( n627 ));
NAND3_X0P5M_A9TL40 U441  (.C ( n628 ) , .Y ( n375 ) , .B ( n359 ));
NAND2_X0P5M_A9TL40 U447  (.B ( n628 ) , .Y ( n369 ));
NOR2XB_X0P5M_A9TL40 U443  (.A ( n628 ) , .Y ( n372 ));
NOR3_X2M_A9TL40 U444  (.B ( n628 ));
NOR3_X0P5M_A9TL40 U417  (.A ( n627 ) , .B ( G33 ) , .Y ( n399 ));
NOR3_X1M_A9TL40 U558  (.A ( n627 ) , .Y ( n428 ));
NOR3_X1A_A9TL40 U553  (.B ( n627 ));
NAND2_X0P5B_A9TL40 U555  (.B ( n627 ) , .A ( n367 ));
INV_X1M_A9TL40 U56  (.A ( n626 ) , .Y ( n625 ));
BUF_X1M_A9TL40 U1  (.A ( n625 ));
INV_X1M_A9TL40 U54  (.A ( n624 ) , .Y ( n623 ));
BUF_X1M_A9TL40 U20  (.A ( n623 ));
INV_X1B_A9TL40 U52  (.A ( n622 ) , .Y ( n621 ));
BUF_X1M_A9TL40 U18  (.A ( n621 ));
INV_X1M_A9TL40 U50  (.A ( n620 ) , .Y ( n619 ));
BUFH_X1M_A9TL40 U16  (.A ( n619 ));
INV_X1B_A9TL40 U48  (.A ( n618 ) , .Y ( n617 ));
BUFH_X1M_A9TL40 U14  (.A ( n617 ));
INV_X0P7B_A9TL40 U46  (.A ( n616 ) , .Y ( n615 ));
BUF_X1M_A9TL40 U12  (.A ( n615 ));
BUF_X1M_A9TL40 U9  (.A ( n614 ));
INV_X1B_A9TL40 U43  (.A ( n613 ) , .Y ( n612 ));
BUFH_X1M_A9TL40 U7  (.A ( n612 ));
INV_X1B_A9TL40 U41  (.A ( n611 ) , .Y ( n610 ));
BUF_X1P2M_A9TL40 U3  (.Y ( n599 ));
BUF_X1M_A9TL40 U5  (.A ( n610 ));
INV_X0P8M_A9TL40 U39  (.A ( n609 ) , .Y ( n608 ));
BUF_X1P2M_A9TL40 U31  (.A ( n608 ));
INV_X0P7B_A9TL40 U37  (.A ( n607 ) , .Y ( n606 ));
BUF_X1P2M_A9TL40 U29  (.A ( n606 ));
INV_X0P8B_A9TL40 U35  (.A ( n605 ) , .Y ( n604 ));
BUFH_X1M_A9TL40 U27  (.A ( n604 ));
INV_X1M_A9TL40 U23  (.A ( n603 ) , .Y ( n602 ));
BUF_X1M_A9TL40 U25  (.A ( n602 ));
DFFRPQ_X0P5M_A9TL40 G29_reg  (.R ( n600 ) , .CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G31_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G32_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G34_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G35_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G36_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G37_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G38_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G39_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G40_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G42_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G43_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G44_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G33_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G41_reg  (.R ( n600 ));
DFFRPQ_X0P5M_A9TL40 G45_reg  (.R ( n600 ) , .Q ( G45 ));
NOR2_X0P5M_A9TL40 U543  (.B ( n256 ) , .Y ( n308 ) , .A ( n414 ));
AOI22_X0P5M_A9TL40 U532  (.B0 ( n256 ) , .Y ( G512 ));
AOI21_X0P5M_A9TL40 U407  (.A1 ( n256 ) , .Y ( n431 ));
OAI211_X0P5M_A9TL40 U456  (.A1 ( n256 ) , .Y ( n392 ));
OR2_X0P7M_A9TL40 U343  (.Y ( n256 ));
AOI21_X0P5M_A9TL40 U433  (.A1 ( n598 ) , .B0 ( n405 ) , .Y ( n411 ));
NAND3_X0P5M_A9TL40 U495  (.A ( n598 ));
AOI22_X0P5M_A9TL40 U532  (.A1 ( n598 ) , .Y ( G512 ));
NAND2_X0P5B_A9TL40 U564  (.B ( n598 ) , .Y ( n430 ));
AOI21_X0P5M_A9TL40 U387  (.A0 ( n598 ) , .B0 ( n325 ) , .Y ( n327 ));
OAI221_X0P5M_A9TL40 U475  (.A1 ( n598 ));
OAI22_X0P5M_A9TL40 U311  (.A0 ( n598 ));
NAND4_X0P5A_A9TL40 U317  (.B ( n598 ) , .C ( G37 ));
NAND2_X0P5B_A9TL40 U357  (.A ( n598 ));
AOI31_X0P5M_A9TL40 U371  (.A1 ( n598 ));
NOR2_X1M_A9TL40 U526  (.Y ( n462 ));
AOI22_X0P5M_A9TL40 U440  (.B1 ( n462 ) , .Y ( n407 ) , .A1 ( n493 ));
AOI21_X0P5M_A9TL40 U403  (.B0 ( n462 ) , .Y ( n324 ));
AO21A1AI2_X0P5M_A9TL40 U467  (.B0 ( n462 ));
NOR3_X0P5M_A9TL40 U303  (.B ( n597 ) , .Y ( n322 ) , .C ( n345 ));
NAND3_X0P5M_A9TL40 U494  (.C ( n597 ));
AOI21_X0P5M_A9TL40 U502  (.A1 ( n597 ) , .B0 ( n294 ) , .Y ( G502 ));
AO21A1AI2_X0P5M_A9TL40 U386  (.A1 ( n597 ) , .Y ( n288 ));
OAI22BB_X0P5M_A9TL40 U392  (.A1 ( n597 ) , .Y ( n393 ));
OAI22_X0P5M_A9TL40 U455  (.A0 ( n597 ) , .Y ( n456 ));
NOR2_X0P5A_A9TL40 U307  (.B ( n597 ));
BUF_X1P2M_A9TL40 U31  (.Y ( n595 ));
NOR2_X0P5M_A9TL40 U565  (.A ( n595 ));
AO21A1AI2_X0P5M_A9TL40 U525  (.A0 ( n595 ) , .Y ( n291 ));
NAND2_X0P5B_A9TL40 U401  (.A ( n595 ));
NAND4_X0P7M_A9TL40 U413  (.A ( n595 ) , .B ( n337 ) , .Y ( n436 ));
NAND2_X0P5B_A9TL40 U414  (.B ( n595 ));
AOI22_X0P5M_A9TL40 U420  (.A0 ( n595 ));
OAI31_X0P7M_A9TL40 U429  (.A0 ( n595 ) , .B0 ( n494 ));
NOR2_X0P7M_A9TL40 U309  (.A ( n595 ));
OAI22_X0P5M_A9TL40 U311  (.B0 ( n595 ));
AOI22_X0P5M_A9TL40 U346  (.A0 ( n595 ));
NOR3_X0P5M_A9TL40 U417  (.C ( n596 ) , .B ( G33 ) , .Y ( n399 ));
OA1B2_X0P5M_A9TL40 U498  (.A0N ( n596 ) , .Y ( n306 ) , .B1 ( n329 ) , .B0 ( n330 ));
NOR2_X0P5M_A9TL40 U527  (.B ( n596 ) , .Y ( n487 ));
NAND2_X0P5B_A9TL40 U480  (.A ( n596 ) , .B ( n448 ) , .Y ( n406 ));
NAND2_X0P5B_A9TL40 U483  (.B ( n596 ) , .Y ( n341 ));
NAND3_X0P5M_A9TL40 U524  (.C ( n596 ));
AOI22_X0P5M_A9TL40 U420  (.B1 ( n596 ));
AO21A1AI2_X0P5M_A9TL40 U467  (.C0 ( n596 ));
OAI31_X0P5M_A9TL40 U469  (.A1 ( n596 ));
OR2_X0P7M_A9TL40 U343  (.B ( n596 ));
OAI21_X0P5M_A9TL40 U355  (.B0 ( n596 ));
BUF_X1P2M_A9TL40 U29  (.Y ( n593 ));
NAND2_X0P5M_A9TL40 U471  (.B ( n593 ) , .Y ( n401 ) , .A ( n488 ));
NAND2_X0P5M_A9TL40 U481  (.B ( n593 ) , .Y ( n400 ));
NOR2_X0P5M_A9TL40 U527  (.A ( n593 ) , .Y ( n487 ));
AO21A1AI2_X0P5M_A9TL40 U567  (.A1 ( n593 ) , .C0 ( n489 ));
OA21A1OI2_X0P5M_A9TL40 U566  (.B0 ( n593 ) , .A1 ( n433 ));
NAND3_X0P5M_A9TL40 U503  (.A ( n593 ) , .Y ( n293 ));
AOI22_X0P5M_A9TL40 U532  (.A0 ( n593 ) , .Y ( G512 ));
NAND2_X1M_A9TL40 U542  (.B ( n593 ));
AOI21_X0P5M_A9TL40 U403  (.A0 ( n593 ) , .Y ( n324 ));
OAI221_X0P5M_A9TL40 U475  (.A0 ( n593 ));
AOI31_X0P5M_A9TL40 U366  (.A0 ( n593 ));
AOI31_X0P5M_A9TL40 U372  (.A0 ( n593 ));
NOR3_X0P5M_A9TL40 U303  (.A ( n594 ) , .Y ( n322 ) , .C ( n345 ));
NAND2_X0P5B_A9TL40 U483  (.A ( n594 ) , .Y ( n341 ));
AOI22_X0P5M_A9TL40 U532  (.B1 ( n594 ) , .Y ( G512 ));
OAI22BB_X0P5M_A9TL40 U392  (.A0 ( n594 ) , .Y ( n393 ));
NOR3_X0P7M_A9TL40 U395  (.C ( n594 ));
OAI22_X0P7M_A9TL40 U430  (.B1 ( n594 ) , .B0 ( n409 ));
AO21A1AI2_X0P5M_A9TL40 U467  (.A1 ( n594 ));
AOI211_X0P7M_A9TL40 U473  (.C0 ( n594 ));
OAI221_X0P5M_A9TL40 U475  (.B0 ( n594 ));
NOR2_X0P5A_A9TL40 U337  (.B ( n594 ));
AOI31_X1M_A9TL40 U369  (.A2 ( n594 ));
BUFH_X1M_A9TL40 U27  (.Y ( n591 ));
NOR2_X0P5M_A9TL40 U331  (.A ( n591 ) , .Y ( n492 ));
NAND3_X0P5M_A9TL40 U524  (.A ( n591 ));
AO21A1AI2_X0P5M_A9TL40 U525  (.C0 ( n591 ) , .Y ( n291 ));
OAI22_X0P5M_A9TL40 U396  (.A0 ( n591 ) , .B0 ( n465 ) , .Y ( n348 ) , .B1 ( n410 ));
NAND2_X0P5B_A9TL40 U414  (.A ( n591 ));
AO21A1AI2_X0P7M_A9TL40 U448  (.C0 ( n591 ) , .B0 ( n452 ));
AO21A1AI2_X0P5M_A9TL40 U467  (.A0 ( n591 ));
OAI31_X0P5M_A9TL40 U469  (.A0 ( n591 ));
AOI211_X0P7M_A9TL40 U473  (.B0 ( n591 ));
OAI31_X1M_A9TL40 U301  (.A0 ( n591 ) , .B0 ( n357 ));
AOI211_X0P5M_A9TL40 U374  (.A0 ( n591 ) , .Y ( G516 ));
NOR3_X0P5M_A9TL40 U496  (.B ( n592 ) , .Y ( n323 ));
AOI22_X0P5M_A9TL40 U440  (.A0 ( n592 ) , .Y ( n407 ) , .A1 ( n493 ));
NOR2_X1B_A9TL40 U438  (.A ( n592 ) , .Y ( n413 ));
OAI22_X0P5M_A9TL40 U499  (.A0 ( n592 ) , .B0 ( n390 ) , .Y ( n307 ) , .B1 ( n429 ));
AOI31_X0P7M_A9TL40 U452  (.B0 ( n592 ) , .A2 ( n391 ));
AOI211_X0P7M_A9TL40 U453  (.B0 ( n592 ) , .Y ( n355 ) , .C0 ( n474 ) , .A1 ( n354 ));
NAND2_X0P5B_A9TL40 U454  (.A ( n592 ));
NOR2_X1B_A9TL40 U323  (.B ( n592 ));
AOI22_X0P5M_A9TL40 U373  (.A0 ( n592 ));
BUF_X1M_A9TL40 U25  (.Y ( n589 ));
OAI31_X2M_A9TL40 U492  (.A0 ( n589 ) , .B0 ( n434 ) , .A1 ( n490 ) , .Y ( G530 ) , .A2 ( n495 ));
AO21A1AI2_X0P5M_A9TL40 U567  (.A0 ( n589 ) , .C0 ( n489 ));
AO21A1AI2_X0P5M_A9TL40 U386  (.C0 ( n589 ) , .Y ( n288 ));
AOI22_X0P5M_A9TL40 U420  (.A1 ( n589 ));
AOI32_X0P5M_A9TL40 U364  (.A0 ( n589 ) , .Y ( G506 ));
AND2_X0P5M_A9TL40 U356  (.B ( n590 ) , .A ( n395 ) , .Y ( n486 ));
NOR2_X0P5M_A9TL40 U360  (.A ( n590 ));
AND4_X0P5M_A9TL40 U478  (.C ( n590 ) , .Y ( G511 ));
AO21A1AI2_X0P5M_A9TL40 U525  (.B0 ( n590 ) , .Y ( n291 ));
NAND4_X0P5A_A9TL40 U474  (.C ( n590 ));
NOR2_X0P7M_A9TL40 U378  (.A ( n590 ));
BUF_X1M_A9TL40 U20  (.Y ( n584 ));
AOI32_X0P7M_A9TL40 U548  (.A1 ( n584 ) , .A0 ( n315 ) , .A2 ( n314 ) , .Y ( n316 ));
AOI22_X0P5M_A9TL40 U536  (.A0 ( n584 ) , .Y ( G515 ));
AOI21_X0P5M_A9TL40 U391  (.A0 ( n584 ) , .A1 ( n363 ));
AO21A1AI2_X0P5M_A9TL40 U458  (.A0 ( n584 ) , .B0 ( n349 ));
AOI31_X1M_A9TL40 U369  (.A0 ( n584 ));
NOR2_X0P5M_A9TL40 U530  (.A ( n585 ) , .Y ( n302 ));
AOI32_X0P7M_A9TL40 U548  (.B1 ( n585 ) , .A0 ( n315 ) , .A2 ( n314 ) , .Y ( n316 ));
OA21_X0P5M_A9TL40 U523  (.A1 ( n585 ) , .Y ( n287 ));
OAI22_X0P5M_A9TL40 U531  (.A1 ( n585 ) , .Y ( G504 ));
OAI211_X0P5M_A9TL40 U537  (.A1 ( n585 ) , .Y ( n299 ));
OAI21_X0P5M_A9TL40 U563  (.A1 ( n585 ) , .Y ( n421 ));
NOR3_X0P7M_A9TL40 U390  (.B ( n585 ));
NAND2_X0P5B_A9TL40 U410  (.A ( n585 ));
OAI22_X0P5M_A9TL40 U466  (.B0 ( n585 ));
NOR2_X0P5A_A9TL40 U337  (.A ( n585 ));
BUF_X1M_A9TL40 U18  (.Y ( n582 ));
NAND2_X0P5M_A9TL40 U535  (.A ( n582 ) , .Y ( n385 ));
NAND3_X0P5M_A9TL40 U486  (.A ( n582 ) , .Y ( n473 ));
AOI211_X1M_A9TL40 U547  (.B0 ( n582 ));
AOI211_X0P5M_A9TL40 U406  (.A0 ( n582 ) , .Y ( n427 ));
NAND2_X0P5B_A9TL40 U418  (.A ( n582 ));
OAI31_X0P5M_A9TL40 U446  (.A0 ( n582 ) , .B0 ( n289 ) , .Y ( n290 ));
NAND4_X0P5A_A9TL40 U474  (.A ( n582 ));
NOR3_X1M_A9TL40 U326  (.A ( n582 ));
AOI31_X0P5M_A9TL40 U354  (.A0 ( n582 ));
NAND2_X3B_A9TL40 U533  (.A ( n583 ) , .Y ( n475 ));
NOR2_X0P5M_A9TL40 U421  (.B ( n583 ) , .Y ( n383 ));
NAND2_X0P5B_A9TL40 U476  (.A ( n583 ) , .Y ( n377 ));
AND4_X0P5M_A9TL40 U478  (.D ( n583 ) , .Y ( G511 ));
NAND3_X0P5M_A9TL40 U490  (.B ( n583 ) , .A ( n419 ));
AO21A1AI2_X0P5M_A9TL40 U501  (.A1 ( n583 ) , .B0 ( n300 ) , .Y ( G513 ));
OA21_X0P5M_A9TL40 U523  (.B0 ( n583 ) , .Y ( n287 ));
OAI22_X0P5M_A9TL40 U531  (.B1 ( n583 ) , .Y ( G504 ));
NAND3B_X0P5M_A9TL40 U404  (.C ( n583 ));
BUFH_X1M_A9TL40 U16  (.Y ( n580 ));
AOI32_X1M_A9TL40 U459  (.A1 ( n580 ) , .A0 ( n441 ) , .A2 ( n312 ) , .Y ( n313 ) , .B0 ( n311 ));
NAND2_X3B_A9TL40 U533  (.B ( n580 ) , .Y ( n475 ));
NOR3_X0P5M_A9TL40 U497  (.A ( n580 ) , .Y ( n303 ) , .C ( n453 ));
OA21_X0P5M_A9TL40 U523  (.A0 ( n580 ) , .Y ( n287 ));
OAI21_X0P5M_A9TL40 U563  (.B0 ( n580 ) , .Y ( n421 ));
OAI22_X0P5M_A9TL40 U402  (.B0 ( n580 ));
NOR3_X0P7M_A9TL40 U415  (.B ( n580 ));
NAND2_X0P5B_A9TL40 U418  (.B ( n580 ));
AOI211_X0P5M_A9TL40 U358  (.A0 ( n580 ));
AOI32_X1M_A9TL40 U459  (.B1 ( n581 ) , .A0 ( n441 ) , .A2 ( n312 ) , .Y ( n313 ) , .B0 ( n311 ));
NAND2_X0P5M_A9TL40 U412  (.A ( n581 ) , .Y ( n297 ));
NOR2_X0P5M_A9TL40 U530  (.B ( n581 ) , .Y ( n302 ));
OA21_X0P5M_A9TL40 U482  (.A0 ( n581 ) , .Y ( n420 ));
OAI22_X0P5M_A9TL40 U493  (.B1 ( n581 ) , .B0 ( n388 ) , .Y ( G547 ) , .A0 ( n389 ));
OAI21_X0P5M_A9TL40 U529  (.A1 ( n581 ) , .Y ( G510 ));
AOI22_X0P5M_A9TL40 U405  (.A1 ( n581 ));
NAND2_X0P5B_A9TL40 U416  (.A ( n581 ) , .Y ( n309 ));
OAI211_X0P5M_A9TL40 U464  (.A1 ( n581 ));
NAND4_X0P5A_A9TL40 U474  (.D ( n581 ));
BUFH_X1M_A9TL40 U14  (.Y ( n578 ));
NOR2_X0P7M_A9TL40 U540  (.A ( n578 ) , .Y ( n332 ));
AO21A1AI2_X0P5M_A9TL40 U501  (.C0 ( n578 ) , .B0 ( n300 ) , .Y ( G513 ));
AOI211_X1M_A9TL40 U547  (.A0 ( n578 ));
OAI21_X0P5M_A9TL40 U563  (.A0 ( n578 ) , .Y ( n421 ));
NAND3_X0P7M_A9TL40 U399  (.A ( n578 ));
NOR3_X0P7M_A9TL40 U415  (.A ( n578 ));
NAND2_X0P5B_A9TL40 U463  (.A ( n578 ));
OAI22_X0P5M_A9TL40 U466  (.A0 ( n578 ));
NAND4XXXB_X1M_A9TL40 U472  (.A ( n578 ));
NAND4_X0P5A_A9TL40 U317  (.A ( n578 ) , .C ( G37 ));
NOR2_X0P5M_A9TL40 U421  (.A ( n579 ) , .Y ( n383 ));
OA21A1OI2_X0P5M_A9TL40 U560  (.A0 ( n579 ) , .Y ( n422 ));
NOR2_X1M_A9TL40 U477  (.B ( n579 ));
OAI21_X0P5M_A9TL40 U400  (.A0 ( n579 ));
OAI211_X0P5M_A9TL40 U464  (.A0 ( n579 ));
NOR3_X1M_A9TL40 U326  (.B ( n579 ));
BUF_X1M_A9TL40 U12  (.Y ( n576 ));
NAND2_X0P5M_A9TL40 U538  (.A ( n576 ) , .B ( G30 ) , .Y ( n298 ));
NOR2_X0P7M_A9TL40 U540  (.B ( n576 ) , .Y ( n332 ));
NAND2_X0P5M_A9TL40 U535  (.B ( n576 ) , .Y ( n385 ));
NOR2_X1M_A9TL40 U477  (.A ( n576 ));
AND4_X0P5M_A9TL40 U478  (.A ( n576 ) , .Y ( G511 ));
OAI22_X0P5M_A9TL40 U531  (.A0 ( n576 ) , .Y ( G504 ));
OAI211_X0P5M_A9TL40 U537  (.B0 ( n576 ) , .Y ( n299 ));
OAI211_X0P5M_A9TL40 U398  (.A0 ( n576 ) , .Y ( n384 ) , .C0 ( n382 ));
NAND2_X0P5B_A9TL40 U416  (.B ( n576 ) , .Y ( n309 ));
NAND2_X0P7B_A9TL40 U470  (.B ( n576 ));
NOR3_X0P5M_A9TL40 U411  (.C ( n577 ) , .B ( n378 ) , .Y ( n362 ));
NOR3_X1M_A9TL40 U546  (.A ( n577 ) , .Y ( n310 ));
OA21_X0P5M_A9TL40 U482  (.A1 ( n577 ) , .Y ( n420 ));
OAI31_X0P5M_A9TL40 U500  (.A2 ( n577 ) , .B0 ( n295 ) , .Y ( n296 ));
NOR3_X0P7M_A9TL40 U415  (.C ( n577 ));
AOI22_X0P5M_A9TL40 U373  (.B1 ( n577 ));
BUFH_X1M_A9TL40 U10  (.Y ( n574 ) , .A ( n573 ));
NAND2_X0P5M_A9TL40 U412  (.B ( n574 ) , .Y ( n297 ));
NOR3_X0P5M_A9TL40 U497  (.B ( n574 ) , .Y ( n303 ) , .C ( n453 ));
NOR3_X1M_A9TL40 U546  (.C ( n574 ) , .Y ( n310 ));
OAI31_X0P5M_A9TL40 U500  (.A1 ( n574 ) , .B0 ( n295 ) , .Y ( n296 ));
OAI21_X0P5M_A9TL40 U529  (.A0 ( n574 ) , .Y ( G510 ));
NAND2_X0P5B_A9TL40 U383  (.B ( n574 ) , .A ( n336 ));
NOR3_X0P7M_A9TL40 U395  (.A ( n574 ));
AOI21_X0P5M_A9TL40 U403  (.A1 ( n574 ) , .Y ( n324 ));
OAI31_X0P7M_A9TL40 U435  (.A0 ( n574 ) , .Y ( n386 ));
OAI31_X0P5M_A9TL40 U446  (.A1 ( n574 ) , .B0 ( n289 ) , .Y ( n290 ));
NAND2_X0P5B_A9TL40 U324  (.A ( n574 ));
AOI211_X0P5M_A9TL40 U358  (.A1 ( n574 ));
NOR2_X0P5M_A9TL40 U488  (.A ( n575 ) , .Y ( n301 ));
NOR2_X1B_A9TL40 U328  (.B ( n575 ));
NOR2_X0P5M_A9TL40 U297  (.A ( n575 ) , .Y ( n387 ));
NAND3_X0P5M_A9TL40 U490  (.C ( n575 ) , .A ( n419 ));
OAI211_X0P5M_A9TL40 U537  (.A0 ( n575 ) , .Y ( n299 ));
AOI22_X0P5M_A9TL40 U539  (.B0 ( n575 ));
AOI22_X0P5M_A9TL40 U388  (.B1 ( n575 ) , .B0 ( G36 ) , .Y ( n342 ) , .A0 ( n467 ));
AOI22_X0P5M_A9TL40 U405  (.B0 ( n575 ));
NAND2_X0P5B_A9TL40 U408  (.B ( n575 ) , .Y ( n466 ));
NOR2_X0P7M_A9TL40 U419  (.B ( n575 ));
OAI22_X0P7M_A9TL40 U436  (.A0 ( n575 ) , .Y ( n408 ));
AOI22_X0P5M_A9TL40 U373  (.B0 ( n575 ));
BUF_X1M_A9TL40 U9  (.Y ( n573 ));
BUFH_X1M_A9TL40 U7  (.Y ( n571 ));
AOI22_X1M_A9TL40 U423  (.A0 ( n571 ) , .B1 ( n497 ) , .A1 ( n498 ));
NOR2_X0P5M_A9TL40 U489  (.A ( n571 ) , .B ( n454 ) , .Y ( n304 ));
NOR2_X1M_A9TL40 U526  (.A ( n571 ));
NAND2_X1M_A9TL40 U542  (.A ( n571 ));
OAI22BB_X0P5M_A9TL40 U392  (.B0N ( n571 ) , .Y ( n393 ));
OAI31_X0P5M_A9TL40 U394  (.A0 ( n571 ) , .B0 ( n333 ) , .Y ( n335 ) , .A2 ( n334 ));
OAI22_X0P5M_A9TL40 U397  (.B0 ( n571 ) , .Y ( n402 ));
OR2_X0P5M_A9TL40 U409  (.B ( n571 ));
AOI22_X0P5M_A9TL40 U420  (.B0 ( n571 ));
NAND2_X0P5B_A9TL40 U462  (.A ( n571 ) , .B ( n326 ));
AOI211_X0P5M_A9TL40 U375  (.A0 ( n571 ));
NOR2_X0P5M_A9TL40 U331  (.B ( n572 ) , .Y ( n492 ));
AOI211_X0P5M_A9TL40 U385  (.A1 ( n572 ) , .B0 ( n484 ) , .C0 ( n483 ));
NAND2_X0P5B_A9TL40 U389  (.A ( n572 ) , .B ( n346 ) , .Y ( n472 ));
NOR3_X0P7M_A9TL40 U390  (.A ( n572 ));
NAND3B_X0P5M_A9TL40 U404  (.B ( n572 ));
NAND4_X0P7M_A9TL40 U413  (.C ( n572 ) , .B ( n337 ) , .Y ( n436 ));
AOI211_X0P7M_A9TL40 U473  (.A0 ( n572 ));
NOR3_X0P5A_A9TL40 U310  (.A ( n572 ) , .Y ( n457 ));
OR2_X0P7M_A9TL40 U343  (.A ( n572 ));
AOI31_X0P5M_A9TL40 U372  (.A1 ( n572 ));
BUF_X1M_A9TL40 U5  (.Y ( n569 ));
AOI22_X1M_A9TL40 U423  (.B0 ( n569 ) , .B1 ( n497 ) , .A1 ( n498 ));
NAND2_X0P5M_A9TL40 U481  (.A ( n569 ) , .Y ( n400 ));
NOR3_X0P5M_A9TL40 U496  (.A ( n569 ) , .Y ( n323 ));
AOI21_X0P5M_A9TL40 U407  (.A0 ( n569 ) , .Y ( n431 ));
NOR2_X0P7M_A9TL40 U419  (.A ( n569 ));
OAI211_X0P5M_A9TL40 U456  (.A0 ( n569 ) , .Y ( n392 ));
OAI211_X0P5M_A9TL40 U460  (.A0 ( n569 ) , .B0 ( n464 ) , .C0 ( n463 ));
OAI221_X0P5M_A9TL40 U475  (.C0 ( n569 ));
NOR2_X1M_A9TL40 U526  (.B ( n570 ));
NOR2_X1B_A9TL40 U328  (.A ( n570 ));
AOI21_X0P7M_A9TL40 U549  (.A1 ( n570 ) , .Y ( n318 ) , .A0 ( n317 ));
AND4_X0P5M_A9TL40 U478  (.B ( n570 ) , .Y ( G511 ));
NAND3_X0P5M_A9TL40 U503  (.C ( n570 ) , .Y ( n293 ));
AO21A1AI2_X0P5M_A9TL40 U525  (.A1 ( n570 ) , .Y ( n291 ));
NAND2_X0P5B_A9TL40 U564  (.A ( n570 ) , .Y ( n430 ));
NAND2_X0P5B_A9TL40 U408  (.A ( n570 ) , .Y ( n466 ));
NAND4_X0P7M_A9TL40 U413  (.D ( n570 ) , .B ( n337 ) , .Y ( n436 ));
AOI211_X0P7M_A9TL40 U431  (.A1 ( n570 ));
NOR2_X1B_A9TL40 U323  (.A ( n570 ));
BUF_X1M_A9TL40 U1  (.Y ( n565 ));
NAND3_X0P5M_A9TL40 U441  (.A ( n565 ) , .Y ( n375 ) , .B ( n359 ));
AOI2XB1_X0P5M_A9TL40 U556  (.B0 ( n565 ) , .A0 ( n439 ) , .Y ( n476 ));
OAI22_X0P5M_A9TL40 U491  (.B0 ( n565 ) , .Y ( G539 ) , .A0 ( n376 ) , .B1 ( n374 ));
NOR3_X1A_A9TL40 U553  (.A ( n565 ));
NOR3_X2M_A9TL40 U444  (.A ( n565 ));
OAI22_X0P5M_A9TL40 U298  (.A0 ( n565 ) , .Y ( n440 ));
AOI32_X0P5M_A9TL40 U364  (.A1 ( n565 ) , .Y ( G506 ));
NOR3_X1M_A9TL40 U558  (.B ( n566 ) , .Y ( n428 ));
NAND2_X0P7M_A9TL40 U437  (.A ( n566 ) , .Y ( n438 ));
AOI32_X0P5M_A9TL40 U364  (.B1 ( n566 ) , .Y ( G506 ));
OA21A1OI2_X0P5M_A9TL40 U566  (.Y ( n434 ) , .A1 ( n433 ));
AO21A1AI2_X0P5M_A9TL40 U567  (.B0 ( n490 ) , .C0 ( n489 ));
NAND3_X0P5M_A9TL40 U524  (.Y ( n490 ));
NOR2_X1B_A9TL40 U461  (.A ( n495 ) , .B ( n347 ) , .Y ( n353 ));
NAND2_X1M_A9TL40 U542  (.Y ( n495 ));
OAI22_X0P5M_A9TL40 U397  (.A1 ( n495 ) , .Y ( n402 ));
AOI31_X0P7M_A9TL40 U424  (.A2 ( n495 ) , .B0 ( n412 ));
OAI31_X0P7M_A9TL40 U429  (.A2 ( n495 ) , .B0 ( n494 ));
NOR2_X1B_A9TL40 U368  (.A ( n495 ));
OAI21_X0P5M_A9TL40 U377  (.A1 ( n495 ) , .Y ( G505 ) , .B0 ( n305 ));
AOI211_X0P5M_A9TL40 U385  (.Y ( n505 ) , .B0 ( n484 ) , .C0 ( n483 ));
OAI211_X0P5M_A9TL40 U426  (.A1 ( n504 ) , .Y ( G549 ) , .A0 ( n398 ) , .B0 ( n397 ) , .C0 ( n396 ));
INV_X0P7B_A9TL40 U294  (.Y ( n504 ));
AOI22_X1M_A9TL40 U423  (.Y ( n503 ) , .B1 ( n497 ) , .A1 ( n498 ));
NAND3_X0P5M_A9TL40 U495  (.Y ( n502 ));
OAI31_X0P7M_A9TL40 U429  (.Y ( n497 ) , .B0 ( n494 ));
AO21A1AI2_X0P5M_A9TL40 U567  (.Y ( n498 ) , .C0 ( n489 ));
AOI22_X0P5M_A9TL40 U440  (.B0 ( n491 ) , .Y ( n407 ) , .A1 ( n493 ));
NAND3_X0P5M_A9TL40 U494  (.B ( n491 ));
NOR3_X1A_A9TL40 U553  (.Y ( n491 ));
AOI21_X0P5M_A9TL40 U293  (.A1 ( n491 ));
AOI22_X0P5M_A9TL40 U365  (.B0 ( n491 ) , .B1 ( G39 ));
AOI31_X0P5M_A9TL40 U371  (.A0 ( n491 ));
NAND2_X0P5M_A9TL40 U361  (.A ( n394 ) , .B ( n482 ) , .Y ( G507 ));
NOR2_X1B_A9TL40 U368  (.B ( n394 ));
NOR2_X0P5M_A9TL40 U565  (.Y ( n470 ));
OA21A1OI2_X0P5M_A9TL40 U566  (.C0 ( n470 ) , .A1 ( n433 ));
INV_X0P6B_A9TL40 U295  (.A ( n470 ) , .Y ( n444 ));
OAI21_X0P5M_A9TL40 U353  (.B0 ( n470 ));
OAI211_X0P5M_A9TL40 U427  (.B0 ( n481 ) , .Y ( G532 ) , .A0 ( G43 ) , .C0 ( n480 ));
AO21B_X0P5M_A9TL40 U457  (.Y ( n469 ) , .A0 ( n468 ));
OAI211_X0P5M_A9TL40 U460  (.Y ( n471 ) , .B0 ( n464 ) , .C0 ( n463 ));
NOR2_X0P5M_A9TL40 U360  (.Y ( n500 ));
NAND3_X0P5M_A9TL40 U495  (.B ( n500 ));
INV_X0P7B_A9TL40 U296  (.A ( n500 ));
NAND3_X0P5M_A9TL40 U503  (.B ( n492 ) , .Y ( n293 ));
AOI21_X0P5M_A9TL40 U407  (.B0 ( n492 ) , .Y ( n431 ));
AOI22_X0P5M_A9TL40 U365  (.A1 ( n492 ) , .B1 ( G39 ));
NAND2_X0P5B_A9TL40 U476  (.B ( n441 ) , .Y ( n377 ));
NOR2_X1M_A9TL40 U477  (.Y ( n441 ));
INV_X0P7B_A9TL40 U327  (.A ( n441 ));
OAI21_X0P5M_A9TL40 U351  (.A0 ( n441 ));
AOI31_X0P5M_A9TL40 U354  (.A1 ( n441 ));
INV_X0P5B_A9TL40 U332  (.Y ( n312 ) , .A ( G31 ));
AOI22_X0P5M_A9TL40 U539  (.A0 ( n312 ));
NAND4XXXB_X1M_A9TL40 U472  (.B ( n312 ));
AOI32_X0P7M_A9TL40 U548  (.B0 ( n313 ) , .A0 ( n315 ) , .A2 ( n314 ) , .Y ( n316 ));
AOI211_X1M_A9TL40 U547  (.Y ( n311 ));
INV_X0P5B_A9TL40 U479  (.A ( n475 ) , .Y ( n381 ));
OA21A1OI2_X0P7M_A9TL40 U450  (.A1 ( n475 ) , .B0 ( n446 ) , .Y ( n344 ));
NAND4XXXB_X1M_A9TL40 U472  (.C ( n475 ));
NOR2_X0P7M_A9TL40 U314  (.A ( n475 ));
NOR2_X0P5A_A9TL40 U379  (.A ( n475 ));
AOI211_X1M_A9TL40 U547  (.A1 ( G31 ));
DFFRPQ_X0P5M_A9TL40 G31_reg  (.Q ( G31 ));
NOR2_X0P5M_A9TL40 U439  (.B ( n375 ) , .Y ( n451 ) , .A ( n366 ));
OAI22_X0P5M_A9TL40 U491  (.A1 ( n375 ) , .Y ( G539 ) , .A0 ( n376 ) , .B1 ( n374 ));
NOR3_X0P5M_A9TL40 U496  (.C ( n359 ) , .Y ( n323 ));
NOR3_X1M_A9TL40 U558  (.C ( n359 ) , .Y ( n428 ));
OAI211_X1M_A9TL40 U550  (.Y ( n359 ) , .A0 ( n338 ) , .A1 ( n319 ) , .B0 ( G46 ));
NOR3_X0P5M_A9TL40 U411  (.A ( n383 ) , .B ( n378 ) , .Y ( n362 ));
OA21_X0P5M_A9TL40 U482  (.B0 ( n383 ) , .Y ( n420 ));
AOI21_X0P5M_A9TL40 U534  (.A0 ( n383 ));
OAI211_X0P5M_A9TL40 U398  (.A1 ( n383 ) , .Y ( n384 ) , .C0 ( n382 ));
OAI22_X0P5M_A9TL40 U397  (.B1 ( n401 ) , .Y ( n402 ));
OAI22_X0P5M_A9TL40 U397  (.A0 ( n488 ) , .Y ( n402 ));
INV_X0P7B_A9TL40 U316  (.A ( n488 ));
NOR2_X1B_A9TL40 U323  (.Y ( n488 ));
AOI31_X0P5M_A9TL40 U348  (.A0 ( n488 ));
INV_X0P5B_A9TL40 U321  (.A ( n297 ) , .Y ( n449 ));
OAI21_X0P5M_A9TL40 U529  (.B0 ( n297 ) , .Y ( G510 ));
OAI211_X0P5M_A9TL40 U537  (.C0 ( n297 ) , .Y ( n299 ));
AOI21_X0P5M_A9TL40 U534  (.A1 ( n449 ));
AOI22_X0P5M_A9TL40 U349  (.B1 ( n449 ));
OAI211_X0P5M_A9TL40 U398  (.B0 ( G34 ) , .Y ( n384 ) , .C0 ( n382 ));
OAI211_X0P5M_A9TL40 U464  (.C0 ( G34 ));
AOI211_X0P5M_A9TL40 U291  (.A0 ( G34 ) , .Y ( G514 ) , .C0 ( n361 ));
DFFRPQ_X0P5M_A9TL40 G34_reg  (.Q ( G34 ));
OA21A1OI2_X0P5M_A9TL40 U560  (.A1 ( n364 ) , .Y ( n422 ));
OAI22_X0P5M_A9TL40 U561  (.A1 ( n364 ) , .B0 ( G42 ) , .Y ( G548 ) , .A0 ( n365 ));
OAI22_X0P5M_A9TL40 U499  (.A1 ( n415 ) , .B0 ( n390 ) , .Y ( n307 ) , .B1 ( n429 ));
AOI31_X0P7M_A9TL40 U452  (.A1 ( n415 ) , .A2 ( n391 ));
NAND2_X0P5B_A9TL40 U324  (.Y ( n415 ));
NAND3_X0P5M_A9TL40 U494  (.A ( n485 ));
AOI211_X0P5M_A9TL40 U385  (.A0 ( n485 ) , .B0 ( n484 ) , .C0 ( n483 ));
OAI31_X0P5M_A9TL40 U469  (.A2 ( n400 ));
AOI31_X0P5M_A9TL40 U371  (.A2 ( n400 ));
NOR2_X0P5M_A9TL40 U488  (.B ( n378 ) , .Y ( n301 ));
OAI21_X0P5M_A9TL40 U400  (.A1 ( n378 ));
OAI31_X0P5M_A9TL40 U449  (.A1 ( n378 ) , .B0 ( n350 ) , .Y ( n356 ) , .A0 ( n351 ));
OAI22_X0P5M_A9TL40 U466  (.A1 ( n378 ));
INV_X0P7B_A9TL40 U330  (.Y ( n378 ));
AOI21_X0P5M_A9TL40 U391  (.B0 ( n362 ) , .A1 ( n363 ));
DFFRPQ_X0P5M_A9TL40 G33_reg  (.Q ( G33 ));
AOI211_X0P7M_A9TL40 U431  (.B0 ( n399 ));
AOI31_X0P5M_A9TL40 U371  (.B0 ( n399 ));
AOI211_X0P5M_A9TL40 U374  (.C0 ( n306 ) , .Y ( G516 ));
OAI31_X1M_A9TL40 U485  (.A2 ( n329 ) , .Y ( n368 ) , .A0 ( n331 ));
AOI211_X0P7M_A9TL40 U473  (.Y ( n329 ));
OAI31_X1M_A9TL40 U485  (.A1 ( n330 ) , .Y ( n368 ) , .A0 ( n331 ));
NOR3_X0P7M_A9TL40 U395  (.Y ( n330 ));
INV_X0P5B_A9TL40 U545  (.A ( G30 ) , .Y ( n321 ));
OAI31_X0P5M_A9TL40 U446  (.A2 ( G30 ) , .B0 ( n289 ) , .Y ( n290 ));
DFFSQN_X0P5M_A9TL40 G30_reg  (.QN ( G30 ));
AOI22_X0P5M_A9TL40 U539  (.B1 ( n298 ));
NAND2XB_X0P5M_A9TL40 U384  (.BN ( n454 ) , .Y ( n445 ));
NAND3_X0P7M_A9TL40 U399  (.Y ( n454 ));
AOI211_X0P7M_A9TL40 U453  (.A0 ( n454 ) , .Y ( n355 ) , .C0 ( n474 ) , .A1 ( n354 ));
OAI22_X0P5M_A9TL40 U455  (.A1 ( n454 ) , .Y ( n456 ));
NAND2XB_X0P5M_A9TL40 U541  (.BN ( n304 ) , .Y ( G509 ));
AOI211_X0P5M_A9TL40 U380  (.A1 ( n304 ) , .Y ( G517 ));
AO21A1AI2_X0P5M_A9TL40 U501  (.A0 ( n301 ) , .B0 ( n300 ) , .Y ( G513 ));
AOI22_X0P5M_A9TL40 U536  (.B0 ( n301 ) , .Y ( G515 ));
AOI211_X0P5M_A9TL40 U374  (.A1 ( n308 ) , .Y ( G516 ));
NOR2_X1B_A9TL40 U328  (.Y ( n414 ));
NAND2_X0P5B_A9TL40 U401  (.B ( n414 ));
AOI31_X0P7M_A9TL40 U424  (.A0 ( n414 ) , .B0 ( n412 ));
INV_X0P7B_A9TL40 U319  (.A ( n414 ));
AOI32_X0P5M_A9TL40 U364  (.A2 ( n323 ) , .Y ( G506 ));
AOI211_X0P5M_A9TL40 U380  (.C0 ( n303 ) , .Y ( G517 ));
NAND2XB_X0P5M_A9TL40 U541  (.A ( n453 ) , .Y ( G509 ));
NAND3B_X0P5M_A9TL40 U404  (.Y ( n453 ));
OAI22_X0P5M_A9TL40 U455  (.B1 ( n453 ) , .Y ( n456 ));
AOI32_X0P5M_A9TL40 U364  (.B0 ( n322 ) , .Y ( G506 ));
NAND2_X0P5M_A9TL40 U552  (.Y ( n345 ) , .B ( G32 ));
NAND2_X0P5M_A9TL40 U447  (.A ( n345 ) , .Y ( n369 ));
NOR3_X1A_A9TL40 U553  (.C ( n345 ));
DFFRPQ_X0P5M_A9TL40 G41_reg  (.Q ( G41 ));
AOI31_X0P5M_A9TL40 U366  (.Y ( n292 ));
DFFSQN_X0P5M_A9TL40 G46_reg  (.D ( n506 ));
INV_X0P6M_A9TL40 U554  (.Y ( n482 ));
NOR2_X1B_A9TL40 U438  (.B ( n482 ) , .Y ( n413 ));
OAI211_X0P5M_A9TL40 U427  (.A1 ( n482 ) , .Y ( G532 ) , .A0 ( G43 ) , .C0 ( n480 ));
OAI22_X0P7M_A9TL40 U436  (.B0 ( n482 ) , .Y ( n408 ));
DFFRPQ_X0P5M_A9TL40 G34_reg  (.D ( G507 ));
NAND3_X0P5M_A9TL40 U490  (.Y ( n358 ) , .A ( n419 ));
OAI31_X1M_A9TL40 U301  (.A2 ( n358 ) , .B0 ( n357 ));
DFFRPQ_X0P5M_A9TL40 G35_reg  (.D ( G508 ));
NAND2_X0P5B_A9TL40 U383  (.Y ( n435 ) , .A ( n336 ));
NOR2_X0P7M_A9TL40 U304  (.B ( n435 ));
NOR3_X1M_A9TL40 U546  (.B ( n321 ) , .Y ( n310 ));
OAI211_X0P5M_A9TL40 U551  (.A1 ( n321 ) , .Y ( n328 ) , .A0 ( n380 ) , .B0 ( n320 ) , .C0 ( n360 ));
AOI22_X0P5M_A9TL40 U405  (.B1 ( n321 ));
AOI211_X1M_A9TL40 U547  (.C0 ( n310 ));
NAND4XXXB_X1M_A9TL40 U472  (.DN ( n310 ));
NAND3_X0P5M_A9TL40 U486  (.B ( n332 ) , .Y ( n473 ));
AOI22_X0P5M_A9TL40 U405  (.A0 ( n332 ));
NAND2_X0P5B_A9TL40 U410  (.B ( n332 ));
NAND4_X0P5A_A9TL40 U474  (.B ( n332 ));
AOI2XB1_X0P5M_A9TL40 U313  (.A0 ( n332 ));
INV_X0P5B_A9TL40 U468  (.A ( n385 ) , .Y ( n423 ));
AOI22_X0P5M_A9TL40 U536  (.B1 ( n385 ) , .Y ( G515 ));
OAI22_X0P5M_A9TL40 U402  (.B1 ( n385 ));
OAI31_X0P7M_A9TL40 U435  (.A2 ( n385 ) , .Y ( n386 ));
AOI211_X0P5M_A9TL40 U358  (.C0 ( n385 ));
NAND3_X0P5M_A9TL40 U486  (.C ( n302 ) , .Y ( n473 ));
OAI22_X0P5M_A9TL40 U531  (.B0 ( n302 ) , .Y ( G504 ));
NAND3_X0P7M_A9TL40 U399  (.C ( n302 ));
INV_X0P7B_A9TL40 U330  (.A ( n302 ));
AOI21_X0P5M_A9TL40 U502  (.A0 ( n487 ) , .B0 ( n294 ) , .Y ( G502 ));
OAI22BB_X0P5M_A9TL40 U392  (.B1N ( n487 ) , .Y ( n393 ));
NOR2_X0P5A_A9TL40 U307  (.A ( n487 ));
NAND2_X0P5B_A9TL40 U324  (.B ( n487 ));
AOI31_X0P5M_A9TL40 U348  (.A1 ( n487 ));
AOI21_X0P5M_A9TL40 U382  (.A0 ( n487 ));
AOI22_X0P5M_A9TL40 U405  (.Y ( n315 ));
NAND4XXXB_X1M_A9TL40 U472  (.Y ( n314 ));
AOI21_X0P7M_A9TL40 U549  (.B0 ( n316 ) , .Y ( n318 ) , .A0 ( n317 ));
NAND3_X0P7M_A9TL40 U399  (.B ( n423 ));
OAI21_X0P5M_A9TL40 U400  (.B0 ( n423 ));
NAND2_X0P5B_A9TL40 U463  (.B ( n423 ));
OAI211_X0P5M_A9TL40 U464  (.B0 ( n423 ));
OAI31_X0P5M_A9TL40 U500  (.A0 ( n381 ) , .B0 ( n295 ) , .Y ( n296 ));
AOI21_X0P5M_A9TL40 U393  (.A0 ( n381 ) , .B0 ( n379 ));
OAI22_X0P5M_A9TL40 U402  (.A0 ( n381 ));
NAND2_X0P7B_A9TL40 U470  (.A ( n381 ));
OAI211_X1M_A9TL40 U550  (.C0 ( n318 ) , .A0 ( n338 ) , .A1 ( n319 ) , .B0 ( G46 ));
AOI22_X0P5M_A9TL40 U420  (.Y ( n317 ));
NAND2_X0P5M_A9TL40 U552  (.A ( n328 ) , .B ( G32 ));
OAI31_X1M_A9TL40 U485  (.B0 ( n328 ) , .Y ( n368 ) , .A0 ( n331 ));
AOI21_X0P5M_A9TL40 U393  (.A1 ( n380 ) , .B0 ( n379 ));
OAI22_X0P5M_A9TL40 U402  (.A1 ( n380 ));
OA21A1OI2_X0P7M_A9TL40 U450  (.A0 ( n380 ) , .B0 ( n446 ) , .Y ( n344 ));
INV_X0P7B_A9TL40 U327  (.Y ( n380 ));
OAI21_X0P5M_A9TL40 U400  (.Y ( n320 ));
OA21A1OI2_X0P5M_A9TL40 U560  (.C0 ( n360 ) , .Y ( n422 ));
NAND2_X0P7B_A9TL40 U470  (.Y ( n360 ));
OAI22_X0P5M_A9TL40 U396  (.A1 ( n347 ) , .B0 ( n465 ) , .Y ( n348 ) , .B1 ( n410 ));
NAND2_X0P5B_A9TL40 U401  (.Y ( n347 ));
INV_X0P7B_A9TL40 U312  (.A ( n347 ));
NAND2XB_X0P5M_A9TL40 U384  (.A ( n353 ) , .Y ( n445 ));
INV_X0P6B_A9TL40 U305  (.A ( n353 ));
AOI22_X0P5M_A9TL40 U381  (.B1 ( n353 ) , .A1 ( G35 ));
DFFRPQ_X0P5M_A9TL40 G32_reg  (.Q ( G32 ));
NAND3_X0P5M_A9TL40 U524  (.B ( n428 ));
INV_X1B_A9TL40 U289  (.A ( n428 ));
OAI22_X0P7M_A9TL40 U436  (.A1 ( n407 ) , .Y ( n408 ));
INV_X0P6M_A9TL40 U554  (.A ( n493 ));
NOR3_X2M_A9TL40 U444  (.Y ( n493 ));
AOI22_X0P5M_A9TL40 U346  (.B0 ( n493 ));
AOI31_X0P5M_A9TL40 U348  (.A2 ( n493 ));
AOI22_X0P5M_A9TL40 U365  (.A0 ( n493 ) , .B1 ( G39 ));
NOR2_X1B_A9TL40 U367  (.B ( n369 ) , .Y ( n432 ) , .A ( n371 ));
INV_X0P6B_A9TL40 U442  (.A ( n369 ) , .Y ( n370 ));
NOR2_X0P5M_A9TL40 U362  (.Y ( n395 ) , .B ( n418 ) , .A ( n499 ));
OAI21_X0P5M_A9TL40 U355  (.A0 ( n395 ));
OA21A1OI2_X0P5M_A9TL40 U566  (.A0 ( n486 ) , .A1 ( n433 ));
AOI211_X0P7M_A9TL40 U431  (.C0 ( n486 ));
AOI22_X0P5M_A9TL40 U346  (.A1 ( n486 ));
AOI31_X0P5M_A9TL40 U348  (.B0 ( n486 ));
NOR2_X0P5M_A9TL40 U297  (.B ( n418 ) , .Y ( n387 ));
NOR2_X0P5M_A9TL40 U360  (.B ( n418 ));
OAI211_X0P7M_A9TL40 U562  (.A1 ( n418 ) , .Y ( G552 ) , .A0 ( G40 ) , .B0 ( n417 ) , .C0 ( n416 ));
OAI22_X0P5M_A9TL40 U561  (.B1 ( n418 ) , .B0 ( G42 ) , .Y ( G548 ) , .A0 ( n365 ));
OAI31_X0P7M_A9TL40 U435  (.A1 ( n418 ) , .Y ( n386 ));
AOI211_X0P5M_A9TL40 U358  (.B0 ( n418 ));
INV_X1B_A9TL40 U289  (.Y ( n418 ));
NAND3_X0P5M_A9TL40 U495  (.C ( n499 ));
NOR3_X0P7M_A9TL40 U395  (.B ( n499 ));
INV_X0P7B_A9TL40 U316  (.Y ( n499 ));
AOI21_X0P5M_A9TL40 U433  (.A0 ( n413 ) , .B0 ( n405 ) , .Y ( n411 ));
AOI31_X0P7M_A9TL40 U424  (.A1 ( n413 ) , .B0 ( n412 ));
INV_X0P7B_A9TL40 U294  (.A ( n413 ));
NAND2_X0P7M_A9TL40 U437  (.B ( n432 ) , .Y ( n438 ));
AOI2XB1_X0P5M_A9TL40 U556  (.A1N ( n432 ) , .A0 ( n439 ) , .Y ( n476 ));
AOI22_X0P5M_A9TL40 U359  (.B0 ( n371 ) , .A0 ( n373 ));
AOI31_X1M_A9TL40 U369  (.Y ( n371 ));
INV_X0P5B_A9TL40 U559  (.A ( n387 ) , .Y ( n426 ));
AOI31_X0P5M_A9TL40 U354  (.A2 ( n387 ));
AOI22_X0P5M_A9TL40 U349  (.A1 ( n451 ));
NAND2XB_X0P5M_A9TL40 U350  (.BN ( n451 ) , .Y ( G518 ));
NAND2_X0P5B_A9TL40 U357  (.B ( n451 ));
AO21A1AI2_X0P7M_A9TL40 U448  (.Y ( n366 ) , .B0 ( n452 ));
INV_X0P6B_A9TL40 U300  (.A ( n366 ));
OA21A1OI2_X0P5M_A9TL40 U560  (.B0 ( n426 ) , .Y ( n422 ));
OAI22_X0P5M_A9TL40 U493  (.A1 ( n426 ) , .B0 ( n388 ) , .Y ( G547 ) , .A0 ( n389 ));
OAI211_X0P7M_A9TL40 U422  (.A1 ( n426 ) , .Y ( G542 ) , .B0 ( n425 ) , .C0 ( n424 ));
AOI211_X0P7M_A9TL40 U431  (.A0 ( n405 ));
OAI21_X0P5M_A9TL40 U355  (.A1 ( n405 ));
NOR2_X1B_A9TL40 U368  (.Y ( n405 ));
OAI22_X0P7M_A9TL40 U430  (.A0 ( n411 ) , .B0 ( n409 ));
NOR2_X0P5M_A9TL40 U565  (.B ( n438 ));
OAI22_X0P5M_A9TL40 U298  (.B0 ( n438 ) , .Y ( n440 ));
AOI31_X0P5M_A9TL40 U348  (.Y ( n489 ));
NAND2_X0P5B_A9TL40 U555  (.Y ( n439 ) , .A ( n367 ));
OAI22_X0P5M_A9TL40 U298  (.A1 ( n439 ) , .Y ( n440 ));
OAI31_X0P5M_A9TL40 U432  (.B0 ( n476 ) , .A1 ( n478 ) , .A0 ( n479 ) , .A2 ( n477 ));
INV_X0P6B_A9TL40 U292  (.A ( n476 ) , .Y ( n460 ));
AOI22_X0P5M_A9TL40 U347  (.A0 ( n476 ));
INV_X0P6B_A9TL40 U290  (.A ( n422 ));
AOI211_X0P5M_A9TL40 U291  (.B0 ( n422 ) , .Y ( G514 ) , .C0 ( n361 ));
DFFRPQ_X0P5M_A9TL40 G40_reg  (.Q ( G40 ));
AOI31_X0P7M_A9TL40 U424  (.Y ( n417 ) , .B0 ( n412 ));
NAND3_X0P5M_A9TL40 U494  (.Y ( n416 ));
AOI31_X0P7M_A9TL40 U428  (.Y ( n433 ));
OAI31_X0P5M_A9TL40 U449  (.A2 ( n377 ) , .B0 ( n350 ) , .Y ( n356 ) , .A0 ( n351 ));
OAI22_X0P5M_A9TL40 U466  (.B1 ( n377 ));
NAND4_X0P5A_A9TL40 U317  (.D ( G511 ) , .C ( G37 ));
DFFRPQ_X0P5M_A9TL40 G38_reg  (.D ( G511 ));
NOR2_X0P7M_A9TL40 U419  (.Y ( n448 ));
INV_X0P7B_A9TL40 U325  (.A ( n448 ));
AOI21_X0P5M_A9TL40 U370  (.A0 ( n448 ));
AOI21_X0P5M_A9TL40 U382  (.A1 ( n448 ));
OAI31_X0P5M_A9TL40 U394  (.A1 ( n406 ) , .B0 ( n333 ) , .Y ( n335 ) , .A2 ( n334 ));
OAI22_X0P7M_A9TL40 U436  (.B1 ( n406 ) , .Y ( n408 ));
OAI211_X0P5M_A9TL40 U456  (.B0 ( n406 ) , .Y ( n392 ));
AOI211_X0P5M_A9TL40 U406  (.B0 ( n420 ) , .Y ( n427 ));
AOI211_X0P5M_A9TL40 U291  (.A1 ( n420 ) , .Y ( G514 ) , .C0 ( n361 ));
AO21A1AI2_X0P5M_A9TL40 U386  (.A0 ( n341 ) , .Y ( n288 ));
OAI211_X0P7M_A9TL40 U445  (.A1 ( n341 ) , .Y ( n343 ) , .B0 ( n340 ));
NOR2XB_X0P5M_A9TL40 U443  (.BN ( n368 ) , .Y ( n372 ));
NOR3_X2M_A9TL40 U444  (.C ( n368 ));
AOI31_X0P7M_A9TL40 U452  (.Y ( n331 ) , .A2 ( n391 ));
INV_X0P6B_A9TL40 U465  (.A ( n473 ));
NOR3_X0P5A_A9TL40 U310  (.C ( n473 ) , .Y ( n457 ));
NOR2_X0P5A_A9TL40 U376  (.A ( n473 ));
AOI21_X0P5M_A9TL40 U534  (.B0 ( n419 ));
AOI211_X0P5M_A9TL40 U406  (.C0 ( n419 ) , .Y ( n427 ));
NOR3_X0P7M_A9TL40 U415  (.Y ( n419 ));
INV_X0P6B_A9TL40 U300  (.Y ( n376 ));
AOI22_X0P5M_A9TL40 U359  (.Y ( n374 ) , .A0 ( n373 ));
AOI31_X0P5M_A9TL40 U354  (.Y ( n388 ));
AOI21_X0P5M_A9TL40 U393  (.Y ( n389 ) , .B0 ( n379 ));
AOI21_X0P5M_A9TL40 U387  (.A1 ( n390 ) , .B0 ( n325 ) , .Y ( n327 ));
NOR3_X0P7M_A9TL40 U390  (.C ( n390 ));
NOR2_X0P7M_A9TL40 U309  (.B ( n390 ));
NOR3_X0P5A_A9TL40 U310  (.B ( n390 ) , .Y ( n457 ));
OAI22_X0P5M_A9TL40 U311  (.A1 ( n390 ));
INV_X0P7B_A9TL40 U319  (.Y ( n390 ));
AOI211_X0P5M_A9TL40 U374  (.B0 ( n307 ) , .Y ( G516 ));
OR2_X0P5M_A9TL40 U409  (.Y ( n429 ));
AOI31_X0P7M_A9TL40 U428  (.A2 ( n429 ));
AOI21_X0P5M_A9TL40 U534  (.Y ( n295 ));
AOI22_X0P5M_A9TL40 U536  (.A1 ( n296 ) , .Y ( G515 ));
AOI22_X0P5M_A9TL40 U539  (.Y ( n300 ));
DFFRPQ_X0P5M_A9TL40 G40_reg  (.D ( G513 ));
OAI31_X0P5M_A9TL40 U469  (.Y ( n294 ));
DFFRPQ_X0P5M_A9TL40 G29_reg  (.D ( G502 ) , .CK ( blif_clk_net ));
OAI31_X0P5M_A9TL40 U469  (.B0 ( n293 ));
DFFSQN_X0P5M_A9TL40 G30_reg  (.D ( n287 ));
AOI31_X0P5M_A9TL40 U366  (.A2 ( n291 ));
DFFRPQ_X0P5M_A9TL40 G37_reg  (.D ( G510 ));
DFFRPQ_X0P5M_A9TL40 G31_reg  (.D ( G504 ));
DFFRPQ_X0P5M_A9TL40 G39_reg  (.D ( G512 ));
DFFRPQ_X0P5M_A9TL40 G42_reg  (.D ( G515 ));
AOI22_X0P5M_A9TL40 U539  (.A1 ( n299 ));
DFFRPQ_X0P5M_A9TL40 G36_reg  (.D ( G509 ));
NAND3B_X0P5M_A9TL40 U404  (.AN ( n338 ));
NAND2_X0P5B_A9TL40 U410  (.Y ( n338 ));
NOR2_X0P7M_A9TL40 U314  (.B ( n338 ));
NAND2_X0P5B_A9TL40 U418  (.Y ( n319 ));
AOI2XB1_X0P5M_A9TL40 U313  (.A1N ( n319 ));
DFFSQN_X0P5M_A9TL40 G46_reg  (.QN ( G46 ));
OAI31_X1M_A9TL40 U301  (.Y ( n367 ) , .B0 ( n357 ));
INV_X0P6B_A9TL40 U363  (.A ( n367 ));
DFFRPQ_X0P5M_A9TL40 G42_reg  (.Q ( G42 ));
AOI21_X0P5M_A9TL40 U391  (.Y ( n365 ) , .A1 ( n363 ));
AOI211_X0P5M_A9TL40 U406  (.A1 ( n421 ) , .Y ( n427 ));
AOI31_X0P7M_A9TL40 U428  (.A1 ( n430 ));
AOI22_X0P5M_A9TL40 U388  (.A1 ( n336 ) , .B0 ( G36 ) , .Y ( n342 ) , .A0 ( n467 ));
INV_X0P7B_A9TL40 U306  (.Y ( n336 ));
OAI211_X0P7M_A9TL40 U445  (.C0 ( n445 ) , .Y ( n343 ) , .B0 ( n340 ));
OAI21_X0P5M_A9TL40 U451  (.B0 ( n445 ) , .Y ( n447 ));
NOR2_X0P7M_A9TL40 U378  (.B ( n445 ));
AO21A1AI2_X0P5M_A9TL40 U386  (.B0 ( n484 ) , .Y ( n288 ));
NOR2_X0P5A_A9TL40 U307  (.Y ( n484 ));
AOI21_X0P5M_A9TL40 U293  (.A0 ( n483 ));
NOR2_X0P7M_A9TL40 U309  (.Y ( n483 ));
AOI211_X0P5M_A9TL40 U375  (.A1 ( n483 ));
AOI22_X0P5M_A9TL40 U373  (.A1 ( n288 ));
OAI22_X0P5M_A9TL40 U311  (.Y ( n325 ));
AOI31_X0P7M_A9TL40 U452  (.A0 ( n327 ) , .A2 ( n391 ));
DFFRPQ_X0P5M_A9TL40 G36_reg  (.Q ( G36 ));
OAI211_X0P7M_A9TL40 U445  (.A0 ( n342 ) , .Y ( n343 ) , .B0 ( n340 ));
NOR3_X0P7M_A9TL40 U390  (.Y ( n467 ));
AO21B_X0P5M_A9TL40 U457  (.A1 ( n467 ) , .A0 ( n468 ));
NAND2_X0P5B_A9TL40 U454  (.B ( n346 ));
INV_X0P7B_A9TL40 U312  (.Y ( n346 ));
OAI21_X0P5M_A9TL40 U377  (.A0 ( n346 ) , .Y ( G505 ) , .B0 ( n305 ));
OA21A1OI2_X0P7M_A9TL40 U450  (.C0 ( n472 ) , .B0 ( n446 ) , .Y ( n344 ));
OAI21_X0P5M_A9TL40 U451  (.A1 ( n472 ) , .Y ( n447 ));
OAI22_X0P5M_A9TL40 U298  (.B1 ( n472 ) , .Y ( n440 ));
NOR2_X0P5A_A9TL40 U376  (.B ( n472 ));
OAI22_X0P5M_A9TL40 U402  (.Y ( n363 ));
AOI211_X0P5M_A9TL40 U375  (.B0 ( n393 ));
AOI21_X0P5M_A9TL40 U382  (.B0 ( n393 ));
OAI22_X0P5M_A9TL40 U466  (.Y ( n379 ));
NAND4_X0P5A_A9TL40 U317  (.Y ( n333 ) , .C ( G37 ));
AO21A1AI2_X0P7M_A9TL40 U448  (.A1 ( n335 ) , .B0 ( n452 ));
NAND4_X0P5A_A9TL40 U474  (.Y ( n334 ));
OR2_X0P5M_A9TL40 U409  (.A ( n465 ));
NAND2_X0P5B_A9TL40 U414  (.Y ( n465 ));
OAI211_X0P5M_A9TL40 U460  (.A1 ( n465 ) , .B0 ( n464 ) , .C0 ( n463 ));
OAI221_X0P5M_A9TL40 U475  (.B1 ( n465 ));
AO21A1AI2_X0P5M_A9TL40 U458  (.C0 ( n348 ) , .B0 ( n349 ));
OAI22_X0P7M_A9TL40 U430  (.A1 ( n410 ) , .B0 ( n409 ));
AOI211_X0P7M_A9TL40 U473  (.A1 ( n410 ));
INV_X0P7B_A9TL40 U325  (.Y ( n410 ));
AOI22_X0P5M_A9TL40 U346  (.B1 ( n402 ));
OAI31_X0P7M_A9TL40 U435  (.B0 ( n384 ) , .Y ( n386 ));
NAND2_X0P5B_A9TL40 U463  (.Y ( n382 ));
OAI22_X0P5M_A9TL40 U311  (.B1 ( n324 ));
OAI211_X0P7M_A9TL40 U422  (.A0 ( n427 ) , .Y ( G542 ) , .B0 ( n425 ) , .C0 ( n424 ));
AOI31_X0P7M_A9TL40 U428  (.A0 ( n431 ));
AOI31_X0P5M_A9TL40 U366  (.A1 ( n431 ));
OAI22_X0P5M_A9TL40 U455  (.B0 ( n466 ) , .Y ( n456 ));
AO21B_X0P5M_A9TL40 U457  (.B0N ( n466 ) , .A0 ( n468 ));
INV_X0P7B_A9TL40 U322  (.A ( n466 ));
AO21A1AI2_X0P7M_A9TL40 U448  (.A0 ( n337 ) , .B0 ( n452 ));
NOR2_X0P5A_A9TL40 U337  (.Y ( n337 ));
OAI31_X1M_A9TL40 U301  (.A1 ( n436 ) , .B0 ( n357 ));
NOR2_X0P7M_A9TL40 U304  (.A ( n436 ));
INV_X0P7B_A9TL40 U315  (.A ( n436 ) , .Y ( n339 ));
NOR3_X1M_A9TL40 U326  (.C ( n309 ));
INV_X0P6B_A9TL40 U290  (.Y ( n425 ));
OAI211_X0P5M_A9TL40 U464  (.Y ( n424 ));
OAI22_X0P7M_A9TL40 U430  (.Y ( n412 ) , .B0 ( n409 ));
DFFRPQ_X0P5M_A9TL40 G29_reg  (.Q ( G29 ) , .CK ( blif_clk_net ));
AOI31_X0P7M_A9TL40 U428  (.B0 ( n496 ));
OAI31_X0P7M_A9TL40 U429  (.A1 ( n496 ) , .B0 ( n494 ));
INV_X0P7B_A9TL40 U296  (.Y ( n496 ));
AOI31_X0P5M_A9TL40 U371  (.Y ( n404 ));
AOI22_X0P5M_A9TL40 U346  (.Y ( n403 ));
AOI211_X0P5M_A9TL40 U375  (.Y ( n398 ));
AOI211_X0P7M_A9TL40 U431  (.Y ( n397 ));
OAI21_X0P5M_A9TL40 U355  (.Y ( n396 ));
DFFRPQ_X0P5M_A9TL40 G43_reg  (.Q ( G43 ));
OAI31_X0P5M_A9TL40 U432  (.Y ( n480 ) , .A1 ( n478 ) , .A0 ( n479 ) , .A2 ( n477 ));
AOI22_X0P5M_A9TL40 U365  (.Y ( n494 ) , .B1 ( G39 ));
AOI21_X0P5M_A9TL40 U293  (.Y ( n409 ));
NOR2_X0P5A_A9TL40 U376  (.Y ( n478 ));
NOR2_X0P7M_A9TL40 U304  (.Y ( n479 ));
AOI22_X0P5M_A9TL40 U347  (.A1 ( n479 ));
NOR2_X0P5A_A9TL40 U379  (.Y ( n477 ));
AOI22_X0P5M_A9TL40 U347  (.B1 ( n450 ));
AOI22_X0P5M_A9TL40 U349  (.B0 ( n450 ));
NAND2_X0P5B_A9TL40 U357  (.Y ( n437 ));
DFFRPQ_X0P5M_A9TL40 G38_reg  (.Q ( G38 ));
AOI31_X0P5M_A9TL40 U354  (.B0 ( n386 ));
AOI21_X0P5M_A9TL40 U293  (.B0 ( n408 ));
AOI22_X0P5M_A9TL40 U359  (.B1 ( n370 ) , .A0 ( n373 ));
AOI22_X0P5M_A9TL40 U359  (.A1 ( n372 ) , .A0 ( n373 ));
AOI31_X1M_A9TL40 U369  (.B0 ( n343 ));
AOI22_X0P5M_A9TL40 U381  (.Y ( n340 ) , .A1 ( G35 ));
AOI22_X0P5M_A9TL40 U373  (.Y ( n289 ));
AOI31_X0P5M_A9TL40 U366  (.B0 ( n290 ));
AOI22_X0P5M_A9TL40 U349  (.A0 ( n452 ));
NOR2_X0P7M_A9TL40 U378  (.Y ( n452 ));
AO21A1AI2_X0P5M_A9TL40 U458  (.Y ( n350 ) , .B0 ( n349 ));
AOI31_X0P5M_A9TL40 U372  (.A2 ( n356 ));
NAND2_X0P5B_A9TL40 U454  (.Y ( n351 ));
OAI21_X0P5M_A9TL40 U451  (.A0 ( n446 ) , .Y ( n447 ));
INV_X0P7B_A9TL40 U306  (.A ( n446 ));
AOI2XB1_X0P5M_A9TL40 U313  (.Y ( n446 ));
AOI31_X1M_A9TL40 U369  (.A1 ( n344 ));
AOI21_X0P5M_A9TL40 U370  (.B0 ( n447 ));
OAI211_X0P5M_A9TL40 U456  (.C0 ( n391 ) , .Y ( n392 ));
NAND2_X0P5B_A9TL40 U462  (.Y ( n391 ) , .B ( n326 ));
AOI31_X0P5M_A9TL40 U372  (.B0 ( n355 ));
INV_X0P6B_A9TL40 U305  (.Y ( n474 ));
NOR2_X0P5A_A9TL40 U379  (.B ( n474 ));
INV_X0P6B_A9TL40 U308  (.Y ( n354 ) , .A ( n352 ));
OAI21_X0P5M_A9TL40 U353  (.A1 ( n456 ));
AOI211_X0P5M_A9TL40 U375  (.C0 ( n392 ));
AO21A1AI2_X0P5M_A9TL40 U458  (.A1 ( n468 ) , .B0 ( n349 ));
AOI2XB1_X0P5M_A9TL40 U313  (.B0 ( n468 ));
NOR3_X1M_A9TL40 U326  (.Y ( n468 ));
OAI21_X0P5M_A9TL40 U351  (.A1 ( n468 ));
AOI21_X0P5M_A9TL40 U370  (.A1 ( n468 ));
INV_X0P6B_A9TL40 U465  (.Y ( n349 ));
AO21A1AI2_X0P5M_A9TL40 U467  (.Y ( n464 ));
OAI221_X0P5M_A9TL40 U475  (.Y ( n463 ));
INV_X0P7B_A9TL40 U322  (.Y ( n326 ));
AOI211_X0P5M_A9TL40 U380  (.A0 ( n326 ) , .Y ( G517 ));
DFFRPQ_X0P5M_A9TL40 G41_reg  (.D ( G514 ));
AOI211_X0P5M_A9TL40 U358  (.Y ( n361 ));
OAI211_X0P5M_A9TL40 U345  (.A1 ( n460 ) , .Y ( G537 ) , .A0 ( n461 ) , .B0 ( n459 ) , .C0 ( n458 ));
NAND2XB_X0P5M_A9TL40 U350  (.A ( n460 ) , .Y ( G518 ));
OAI211_X0P5M_A9TL40 U344  (.A1 ( n444 ) , .Y ( G535 ) , .A0 ( G44 ) , .B0 ( n443 ) , .C0 ( n442 ));
OAI21_X0P5M_A9TL40 U351  (.B0 ( n440 ));
AOI31_X0P5M_A9TL40 U372  (.Y ( n357 ));
NOR2_X0P7M_A9TL40 U314  (.Y ( n352 ));
AOI22_X0P5M_A9TL40 U381  (.B0 ( n352 ) , .A1 ( G35 ));
OAI21_X0P5M_A9TL40 U353  (.A0 ( n457 ));
AOI211_X0P5M_A9TL40 U380  (.B0 ( n457 ) , .Y ( G517 ));
AOI22_X0P5M_A9TL40 U381  (.A0 ( n339 ) , .A1 ( G35 ));
AOI22_X0P5M_A9TL40 U347  (.B0 ( G37 ));
DFFRPQ_X0P5M_A9TL40 G37_reg  (.Q ( G37 ));
DFFRPQ_X0P5M_A9TL40 G44_reg  (.Q ( G44 ));
AOI22_X0P5M_A9TL40 U347  (.Y ( n443 ));
OAI21_X0P5M_A9TL40 U351  (.Y ( n442 ));
AOI21_X0P5M_A9TL40 U370  (.Y ( n461 ));
AOI22_X0P5M_A9TL40 U349  (.Y ( n459 ));
OAI21_X0P5M_A9TL40 U353  (.Y ( n458 ));
DFFRPQ_X0P5M_A9TL40 G45_reg  (.D ( G518 ) , .Q ( G45 ));
INV_X0P6B_A9TL40 U363  (.Y ( n373 ));
DFFRPQ_X0P5M_A9TL40 G33_reg  (.D ( G506 ));
DFFRPQ_X0P5M_A9TL40 G39_reg  (.Q ( G39 ));
DFFRPQ_X0P5M_A9TL40 G43_reg  (.D ( G516 ));
DFFRPQ_X0P5M_A9TL40 G32_reg  (.D ( G505 ));
AOI21_X0P5M_A9TL40 U382  (.Y ( n305 ));
DFFRPQ_X0P5M_A9TL40 G44_reg  (.D ( G517 ));
DFFRPQ_X0P5M_A9TL40 G35_reg  (.Q ( G35 ));
DFFRPQ_X0P5M_A9TL40 G31_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G32_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G34_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G35_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G36_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G37_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G38_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G39_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G40_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G42_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G43_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G44_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G33_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G41_reg  (.CK ( blif_clk_net ));
DFFRPQ_X0P5M_A9TL40 G45_reg  (.CK ( blif_clk_net ) , .Q ( G45 ));
DFFSQN_X0P5M_A9TL40 G46_reg  (.CK ( blif_clk_net ));
DFFSQN_X0P5M_A9TL40 G30_reg  (.CK ( blif_clk_net ));
endmodule
